/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:24:21 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__21,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire  inst_cellmath__46;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__68,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire N493,N494,N548,N549,N550,N551,N585 
	,N594,N595,N623,N624,N625,N626,N627,N628 
	,N629,N630,N631,N632,N633,N634,N635,N636 
	,N637,N638,N639,N640,N641,N642,N643,N644 
	,N645,N646,N647,N648,N649,N650,N651,N652 
	,N677,N678,N679,N680,N681,N682,N683,N684 
	,N685,N686,N687,N688,N689,N690,N691,N692 
	,N693,N694,N695,N696,N697,N698,N699,N700 
	,N701,N702,N703,N704,N705,N706,N707,N708 
	,N709,N710,N711,N712,N713,N717,N718,N719 
	,N720,N721,N722,N723,N724,N725,N726,N727 
	,N728,N729,N730,N731,N732,N733,N734,N735 
	,N736,N737,N738,N739,N741,N742,N743,N744 
	,N745,N746,N747,N748,N749,N750,N751,N752 
	,N753,N754,N755,N756,N757,N758,N759,N760 
	,N761,N762,N763,N3933,N3934,N3935,N3936,N3937 
	,N3938,N3939,N3940,N3944,N3945,N3946,N3947,N3948 
	,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3957 
	,N3958,N3959,N3960,N3961,N3962,N3963,N3965,N3966 
	,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975 
	,N3976,N3977,N3978,N3979,N3980,N3983,N3984,N3985 
	,N3986,N3987,N3988,N3989,N3990,N3992,N3993,N3994 
	,N3995,N3996,N3998,N3999,N4000,N4001,N4002,N4004 
	,N4005,N4006,N4007,N4008,N4009,N4011,N4012,N4013 
	,N4014,N4015,N4016,N4017,N4018,N4021,N4022,N4023 
	,N4024,N4025,N4027,N4028,N4029,N4030,N4031,N4032 
	,N4033,N4036,N4037,N4038,N4039,N4040,N4041,N4042 
	,N4043,N4045,N4046,N4047,N4048,N4049,N4051,N4052 
	,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4062 
	,N4063,N4064,N4065,N4066,N4067,N4069,N4070,N4071 
	,N4072,N4073,N4075,N4076,N4077,N4078,N4079,N4080 
	,N4081,N4082,N4083,N4085,N4086,N4088,N4089,N4090 
	,N4091,N4092,N4093,N4095,N4096,N4097,N4098,N4099 
	,N4100,N4101,N4102,N4103,N4104,N4105,N4107,N4109 
	,N4110,N4112,N4113,N4114,N4115,N4116,N4117,N4118 
	,N4119,N4120,N4121,N4123,N4124,N4126,N4127,N4128 
	,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136 
	,N4137,N4138,N4139,N4141,N4142,N4145,N4146,N4147 
	,N4148,N4149,N4150,N4151,N4154,N4155,N4156,N4157 
	,N4158,N4160,N4161,N4162,N4163,N4165,N4166,N4167 
	,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176 
	,N4177,N4178,N4179,N4181,N4182,N4183,N4184,N4185 
	,N4186,N4187,N4190,N4191,N4192,N4193,N4194,N4195 
	,N4197,N4198,N4199,N4200,N4201,N4202,N4204,N4205 
	,N4206,N4207,N4208,N4209,N4210,N4211,N4213,N4214 
	,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222 
	,N4223,N4224,N4225,N4226,N4227,N4229,N4230,N4231 
	,N4232,N4234,N4235,N4236,N4237,N4238,N4239,N4241 
	,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249 
	,N4250,N4252,N4253,N4254,N4255,N4256,N4257,N4258 
	,N4260,N4261,N4262,N4263,N4264,N4266,N4268,N4270 
	,N4271,N4272,N4273,N4274,N4275,N4276,N4279,N4280 
	,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4290 
	,N4291,N4292,N4293,N4294,N4295,N4297,N4298,N4299 
	,N4300,N4301,N4302,N4304,N4305,N4306,N4308,N4309 
	,N4310,N4311,N4312,N4313,N4314,N4316,N4317,N4318 
	,N4319,N4320,N4322,N4323,N4324,N4325,N4326,N4329 
	,N4330,N4331,N4333,N4334,N4335,N4336,N4337,N4338 
	,N4339,N4341,N4343,N4344,N4345,N4346,N4347,N4348 
	,N4349,N4350,N4351,N4352,N4353,N4355,N4356,N4359 
	,N4360,N4361,N4363,N4364,N4365,N4366,N4367,N4368 
	,N4369,N4371,N4372,N4373,N4376,N4377,N4378,N4379 
	,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387 
	,N4388,N4389,N4391,N4392,N4393,N4394,N4395,N4396 
	,N4397,N4398,N4399,N4400,N4402,N4403,N4404,N4406 
	,N4407,N4409,N4410,N4411,N4413,N4414,N4415,N4417 
	,N4418,N4419,N4420,N4421,N4422,N4423,N4425,N4426 
	,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434 
	,N4435,N4437,N4438,N4439,N4440,N4441,N4442,N4443 
	,N4444,N4445,N4446,N4447,N4448,N4449,N4451,N4452 
	,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460 
	,N4463,N4464,N4466,N4467,N4468,N4470,N4471,N4472 
	,N4473,N4474,N4476,N4478,N4479,N4480,N4481,N4482 
	,N4484,N4485,N4486,N4488,N4489,N4490,N4493,N4494 
	,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4503 
	,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511 
	,N4513,N4514,N4515,N4516,N4518,N4519,N4520,N4521 
	,N4522,N4524,N4525,N4526,N4527,N4529,N4530,N4532 
	,N4533,N4534,N4535,N4536,N4537,N4538,N4540,N4541 
	,N4542,N4543,N4545,N4546,N4547,N4548,N4549,N4550 
	,N4551,N4552,N4554,N4555,N4556,N4557,N4559,N4560 
	,N4562,N4563,N4565,N4566,N4567,N4568,N4569,N4571 
	,N4573,N4574,N4575,N4576,N4577,N4579,N4580,N4581 
	,N4582,N4584,N4586,N4587,N4588,N4590,N4591,N4592 
	,N4594,N4595,N4596,N4597,N4599,N4600,N4601,N4602 
	,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4611 
	,N4612,N4613,N4614,N4615,N4617,N4618,N4619,N4621 
	,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629 
	,N4630,N4631,N4632,N4634,N4635,N4636,N4638,N4639 
	,N4640,N4641,N4643,N4645,N4647,N4648,N4649,N4650 
	,N4651,N4652,N4653,N4654,N4655,N4657,N4658,N5364 
	,N5371,N5372,N5373,N5376,N5379,N5385,N5402,N5403 
	,N5404,N5405,N5406,N5408,N5409,N5411,N5413,N5414 
	,N5415,N5416,N5417,N5419,N5422,N5423,N5424,N5425 
	,N5427,N5428,N5430,N5431,N5433,N5434,N5435,N5436 
	,N5438,N5440,N5441,N5442,N5443,N5444,N5446,N5447 
	,N5449,N5450,N5451,N5452,N5453,N5455,N5456,N5458 
	,N5459,N5461,N5462,N5463,N5464,N5465,N5467,N5470 
	,N5471,N5472,N5473,N5474,N5476,N5478,N5479,N5481 
	,N5482,N5483,N5485,N5486,N5487,N5489,N5490,N5491 
	,N5493,N5494,N5497,N5498,N5499,N5500,N5501,N5503 
	,N5504,N5505,N5507,N5509,N5510,N5511,N5512,N5513 
	,N5515,N5518,N5519,N5520,N5521,N5523,N5525,N5526 
	,N5527,N5528,N5530,N5531,N5532,N5534,N5535,N5537 
	,N5538,N5539,N5540,N5542,N5545,N5546,N5547,N5549 
	,N5550,N5552,N5553,N5554,N5556,N5557,N5558,N5560 
	,N5562,N5563,N5564,N5565,N5566,N5568,N5569,N5571 
	,N5573,N5574,N5576,N5577,N5578,N5580,N5581,N5583 
	,N5584,N5585,N5586,N5587,N5591,N5592,N5593,N5594 
	,N5595,N5597,N5598,N5599,N5601,N5602,N5604,N5605 
	,N5606,N5608,N5610,N5611,N5612,N5613,N5615,N5616 
	,N5817,N5876,N5877,N5878,N5879,N5880,N5881,N5882 
	,N5883,N5884,N5885,N5886,N5887,N5888,N5890,N5891 
	,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899 
	,N5900,N5901,N5903,N5904,N5905,N5906,N5907,N5908 
	,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5917 
	,N5918,N5920,N5921,N5922,N5923,N5924,N5925,N5926 
	,N5927,N5928,N5929,N5931,N5933,N5934,N5935,N5936 
	,N5937,N5938,N5939,N5940,N5941,N5942,N5944,N5945 
	,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954 
	,N5955,N5957,N5958,N5959,N5960,N5961,N5962,N5963 
	,N5964,N5965,N5966,N5967,N5968,N5970,N5971,N5972 
	,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980 
	,N5981,N5983,N5984,N5985,N5986,N5988,N5989,N5990 
	,N5991,N5992,N5993,N5994,N5995,N5996,N5997,N5998 
	,N5999,N6000,N6002,N6003,N6004,N6005,N6006,N6007 
	,N6008,N6009,N6010,N6011,N6012,N6013,N6015,N6016 
	,N6017,N6019,N6020,N6021,N6022,N6023,N6024,N6025 
	,N6026,N6027,N6028,N6030,N6031,N6033,N6034,N6035 
	,N6036,N6037,N6038,N6039,N6040,N6042,N6043,N6044 
	,N6045,N6046,N6047,N6048,N6049,N6050,N6051,N6052 
	,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060 
	,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068 
	,N6069,N6070,N6071,N6072,N6074,N6075,N6076,N6077 
	,N6078,N6079,N6081,N6082,N6083,N6085,N6086,N6087 
	,N6088,N6090,N6091,N6092,N6093,N6094,N6095,N6096 
	,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6106 
	,N6107,N6108,N6110,N6111,N6112,N6113,N6114,N6115 
	,N6116,N6117,N6119,N6120,N6121,N6122,N6123,N6124 
	,N6125,N6126,N6127,N6128,N6129,N6131,N6132,N6133 
	,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141 
	,N6142,N6144,N6145,N6146,N6147,N6148,N6149,N6150 
	,N6151,N6152,N6153,N6154,N6155,N6156,N6159,N6160 
	,N6161,N6162,N6163,N6164,N6166,N6167,N6168,N6171 
	,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179 
	,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188 
	,N6189,N6190,N6191,N6192,N6193,N6195,N6197,N6198 
	,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206 
	,N6207,N6209,N6210,N6211,N6212,N6213,N6214,N6215 
	,N6216,N6217,N6218,N6219,N6220,N6221,N6223,N6224 
	,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232 
	,N6234,N6235,N6237,N6238,N6239,N6240,N6241,N6242 
	,N6243,N6244,N6245,N6246,N6248,N6250,N6251,N6252 
	,N6253,N6254,N6255,N6256,N6258,N6259,N6260,N6261 
	,N6262,N6264,N6265,N6266,N6267,N6268,N6269,N6270 
	,N6272,N6273,N6274,N6275,N6276,N6277,N6278,N6279 
	,N6280,N6281,N6282,N6283,N6285,N6286,N6287,N6288 
	,N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296 
	,N6297,N6298,N6299,N6301,N6302,N6303,N6304,N6305 
	,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6314 
	,N6315,N6316,N6317,N6318,N6320,N6321,N6322,N6324 
	,N6325,N6326,N6328,N6329,N6330,N6331,N6332,N6333 
	,N6334,N6335,N6337,N6339,N6340,N6341,N6342,N6343 
	,N6344,N6345,N6346,N6348,N6349,N6350,N6351,N6352 
	,N6354,N6355,N6356,N6357,N6358,N6359,N6360,N6361 
	,N6362,N6363,N6365,N6366,N6367,N6368,N6369,N6370 
	,N6371,N6372,N6373,N6374,N6376,N6377,N6378,N6379 
	,N6380,N6381,N6382,N6383,N6385,N6386,N6387,N6388 
	,N6389,N6391,N6392,N6393,N6394,N6395,N6396,N6398 
	,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6407 
	,N6408,N6410,N6411,N6412,N6413,N6414,N6415,N6416 
	,N6417,N6418,N6420,N6421,N6422,N6423,N6424,N6425 
	,N6426,N6427,N6428,N6429,N6431,N6432,N6433,N6434 
	,N6435,N6436,N6437,N6438,N6439,N6440,N6441,N6442 
	,N6443,N6444,N6446,N6447,N6448,N6449,N6450,N6451 
	,N6452,N6453,N6454,N6455,N6456,N6458,N6459,N6460 
	,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6469 
	,N6470,N6471,N6472,N6474,N6475,N6476,N6477,N6478 
	,N6479,N6480,N6481,N6483,N6484,N6485,N6486,N6487 
	,N6488,N6489,N6490,N6491,N6492,N6493,N6494,N6495 
	,N6496,N6499,N6501,N6502,N6503,N6504,N6505,N6506 
	,N6507,N6508,N6509,N6510,N6511,N6513,N6514,N6515 
	,N6516,N6517,N6518,N6519,N6520,N6521,N6522,N6523 
	,N6525,N6526,N6527,N6528,N6529,N6530,N6531,N6532 
	,N6533,N6534,N6536,N6537,N6538,N6539,N6541,N6542 
	,N6543,N6544,N6545,N6546,N6547,N6548,N6550,N6552 
	,N6553,N6554,N6555,N6556,N6558,N6559,N6560,N6561 
	,N6562,N6564,N6565,N6566,N6567,N6568,N6569,N6570 
	,N6571,N6573,N6574,N6575,N6576,N6577,N6578,N6579 
	,N6580,N6581,N6582,N7286,N7287,N7288,N7289,N7290 
	,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7299 
	,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307 
	,N7308,N7310,N7311,N7312,N7313,N7314,N7315,N7316 
	,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324 
	,N7325,N7326,N7327,N7328,N7329,N7330,N7331,N7332 
	,N7333,N7335,N7336,N7337,N7338,N7339,N7340,N7341 
	,N7342,N7343,N7344,N7345,N7346,N7347,N7348,N7349 
	,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7358 
	,N7359,N7362,N7363,N7364,N7365,N7366,N7368,N7369 
	,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377 
	,N7378,N7379,N7380,N7381,N7383,N7385,N7386,N7387 
	,N7388,N7390,N7391,N7392,N7393,N7394,N7395,N7396 
	,N7397,N7398,N7399,N7400,N7402,N7403,N7404,N7405 
	,N7406,N7407,N7408,N7409,N7410,N7411,N7413,N7414 
	,N7416,N7417,N7419,N7420,N7421,N7422,N7424,N7425 
	,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7434 
	,N7435,N7436,N7437,N7438,N7440,N7442,N7443,N7444 
	,N7447,N7448,N7451,N7452,N7454,N7455,N7456,N7457 
	,N7458,N7459,N7460,N7462,N7463,N7464,N7465,N7466 
	,N7467,N7468,N7469,N7470,N7471,N7472,N7473,N7476 
	,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485 
	,N7486,N7487,N7488,N7489,N7490,N7491,N7492,N7493 
	,N7494,N7495,N7496,N7497,N7498,N7499,N7500,N7502 
	,N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7511 
	,N7512,N7513,N7514,N7515,N7516,N7517,N7518,N7519 
	,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527 
	,N7528,N7531,N7532,N7533,N7534,N7535,N7537,N7538 
	,N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546 
	,N7547,N7549,N7550,N7551,N7552,N7553,N7554,N7555 
	,N7556,N7557,N7559,N7560,N7561,N7562,N7563,N7564 
	,N7565,N7566,N7567,N7568,N7569,N7570,N7571,N7572 
	,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580 
	,N7581,N7582,N7584,N7585,N7586,N7587,N7588,N7590 
	,N7591,N7592,N7594,N7595,N7596,N7597,N7598,N7599 
	,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607 
	,N7608,N7609,N7610,N7611,N7612,N7613,N7614,N7615 
	,N7616,N7617,N7619,N7620,N7622,N7623,N7624,N7625 
	,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633 
	,N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641 
	,N7643,N7644,N7645,N7646,N7647,N7648,N7650,N7652 
	,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661 
	,N7663,N7665,N7666,N7667,N7668,N7669,N7670,N7671 
	,N7672,N7674,N7676,N7678,N7679,N7680,N7681,N7682 
	,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690 
	,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698 
	,N7699,N7701,N7702,N7703,N7704,N7705,N7706,N7707 
	,N7708,N7709,N7710,N7712,N7713,N7714,N7715,N7716 
	,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7725 
	,N7726,N7727,N7728,N7729,N7730,N7731,N7733,N7734 
	,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742 
	,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751 
	,N7752,N7753,N7754,N7756,N7757,N7758,N7759,N7760 
	,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768 
	,N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776 
	,N7777,N7779,N7780,N7781,N7782,N7784,N7785,N7786 
	,N7787,N7788,N7789,N7790,N7791,N7792,N7793,N7795 
	,N7796,N7797,N7798,N7799,N7800,N7801,N7804,N7805 
	,N7806,N7807,N7808,N7810,N7811,N7812,N7813,N7814 
	,N7816,N7817,N7818,N7819,N7820,N7822,N7823,N7824 
	,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832 
	,N7833,N7835,N7836,N7837,N7838,N7840,N7841,N7842 
	,N7843,N7844,N7845,N7847,N7849,N7850,N7851,N7852 
	,N7853,N7854,N7855,N7857,N7858,N7859,N7860,N7861 
	,N7863,N7865,N7866,N7867,N7868,N7869,N7870,N7872 
	,N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881 
	,N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889 
	,N7890,N7891,N7892,N7893,N7895,N7896,N7897,N7899 
	,N7900,N7902,N7903,N7904,N7905,N7906,N7907,N7908 
	,N7909,N7910,N7911,N7912,N7914,N7915,N7916,N7917 
	,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925 
	,N7926,N7927,N7929,N7931,N7932,N7933,N7934,N7935 
	,N7936,N7938,N7939,N7940,N8579,N8580,N8581,N8582 
	,N8583,N8585,N8586,N8587,N8588,N8589,N8590,N8591 
	,N8592,N8593,N8594,N8595,N8596,N8597,N8598,N8599 
	,N8600,N8601,N8602,N8603,N8605,N8606,N8607,N8608 
	,N8609,N8610,N8611,N8613,N8615,N8616,N8617,N8618 
	,N8619,N8620,N8621,N8622,N8623,N8624,N8625,N8626 
	,N8627,N8629,N8630,N8631,N8632,N8634,N8635,N8637 
	,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645 
	,N8646,N8647,N8648,N8649,N8650,N8651,N8653,N8654 
	,N8655,N8656,N8657,N8658,N8659,N8660,N8661,N8662 
	,N8663,N8664,N8665,N8666,N8667,N8668,N8670,N8671 
	,N8672,N8673,N8674,N8675,N8676,N8678,N8679,N8680 
	,N8681,N8682,N8685,N8686,N8687,N8688,N8689,N8690 
	,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698 
	,N8699,N8700,N8701,N8703,N8704,N8705,N8706,N8707 
	,N8708,N8710,N8711,N8712,N8713,N8714,N8715,N8716 
	,N8717,N8719,N8721,N8722,N8723,N8724,N8725,N8726 
	,N8727,N8728,N8730,N8731,N8732,N8733,N8734,N8735 
	,N8736,N8739,N8740,N8741,N8742,N8743,N8744,N8745 
	,N8746,N8747,N8748,N8749,N8750,N8751,N8752,N8753 
	,N8754,N8756,N8757,N8758,N8760,N8762,N8763,N8764 
	,N8765,N8766,N8767,N8768,N8769,N8770,N8771,N8772 
	,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780 
	,N8781,N8782,N8783,N8784,N8785,N8787,N8788,N8789 
	,N8790,N8791,N8792,N8793,N8795,N8796,N8797,N8798 
	,N8799,N8800,N8802,N8803,N8804,N8805,N8806,N8807 
	,N8808,N8809,N8810,N8811,N8812,N8813,N8814,N8816 
	,N8817,N8818,N8820,N8822,N8823,N8824,N8825,N8826 
	,N8827,N8828,N8829,N8831,N8832,N8833,N8834,N8835 
	,N8836,N8837,N8838,N8839,N8840,N8841,N8842,N8844 
	,N8845,N8846,N8847,N8849,N8850,N8851,N8852,N8853 
	,N8854,N8855,N8856,N8857,N8858,N8859,N8860,N8862 
	,N8863,N8864,N8865,N8866,N8867,N8868,N8869,N8870 
	,N8871,N8872,N8873,N8875,N8876,N8877,N8880,N8881 
	,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8889 
	,N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897 
	,N8898,N8899,N8900,N8901,N8902,N8904,N8905,N8906 
	,N8907,N8908,N8910,N8911,N8912,N8913,N8914,N8915 
	,N8916,N8917,N8918,N8919,N8920,N8921,N8922,N8923 
	,N8924,N8925,N8926,N8927,N8928,N8929,N8930,N8931 
	,N8932,N8933,N8934,N8935,N8936,N8937,N8938,N8940 
	,N8941,N8942,N8943,N8945,N8946,N8947,N8948,N8949 
	,N8951,N8952,N8953,N8954,N8955,N8956,N8957,N8958 
	,N8959,N8960,N8961,N8962,N8963,N8965,N8966,N8967 
	,N8969,N8970,N8972,N8973,N8974,N8975,N8976,N8977 
	,N8978,N8979,N8980,N8981,N8982,N8983,N8984,N8985 
	,N8986,N8987,N8988,N8989,N8990,N8991,N8992,N8994 
	,N8995,N8996,N8997,N8998,N8999,N9000,N9001,N9002 
	,N9003,N9004,N9005,N9006,N9007,N9008,N9010,N9011 
	,N9012,N9013,N9014,N9015,N9016,N9017,N9018,N9019 
	,N9020,N9021,N9022,N9023,N9024,N9026,N9027,N9028 
	,N9030,N9031,N9032,N9033,N9034,N9035,N9036,N9037 
	,N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045 
	,N9046,N9047,N9048,N9049,N9050,N9051,N9052,N9054 
	,N9055,N9056,N9057,N9058,N9059,N9060,N9062,N9063 
	,N9064,N9065,N9066,N9067,N9068,N9069,N9071,N9072 
	,N9073,N9074,N9075,N9076,N9077,N9078,N9079,N9080 
	,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9089 
	,N9090,N9091,N9092,N9093,N9094,N9096,N9098,N9099 
	,N9100,N9101,N9102,N9103,N9104,N9105,N9106,N9107 
	,N9108,N9109,N9110,N9111,N9112,N9113,N9114,N9115 
	,N9116,N9118,N9119,N9120,N9121,N9122,N9123,N9124 
	,N9126,N9128,N9129,N9130,N9131,N9132,N9133,N9134 
	,N9135,N9136,N9137,N9138,N9139,N9140,N9141,N9143 
	,N9144,N9145,N9146,N9147,N9148,N9149,N9150,N9151 
	,N9152,N9153,N9155,N9156,N9157,N9158,N9159,N9162 
	,N9163,N9164,N9165,N9166,N9168,N9169,N9171,N9172 
	,N9173,N9174,N9175,N9176,N9177,N9178,N9179,N9180 
	,N9181,N9182,N9183,N9185,N9186,N9187,N9188,N9189 
	,N9190,N9192,N9194,N9195,N9196,N9197,N9198,N9199 
	,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207 
	,N9208,N9209,N9210,N9212,N9213,N9214,N9215,N9216 
	,N9217,N9218,N9220,N9221,N9222,N9223,N9224,N9225 
	,N9226,N9227,N9228,N9229,N9230,N9231,N9233,N9234 
	,N9235,N9236,N9237,N9238,N9239,N9240,N9241,N9242 
	,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250 
	,N9251,N9253,N9254,N9255,N9256,N9257,N9258,N9259 
	,N9262,N9263,N9264,N9265,N9266,N9267,N9268,N9269 
	,N9270,N9271,N9272,N9273,N9274,N9275,N9276,N9277 
	,N9278,N9280,N9281,N9282,N9283,N9284,N9285,N9286 
	,N9288,N9289,N9290,N9291,N9292,N9293,N9294,N9295 
	,N9296,N9297,N9298,N9299,N9301,N9302,N9303,N9304 
	,N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312 
	,N9313,N9314,N9315,N9316,N9318,N9319,N9320,N9321 
	,N9322,N9323,N9324,N9325,N9326,N9329,N9330,N9331 
	,N9332,N9333,N9334,N9335,N9336,N9337,N9338,N9339 
	,N9340,N9341,N9342,N9343,N9344,N9346,N9347,N9348 
	,N9349,N9350,N9352,N9353,N9355,N9356,N9357,N9358 
	,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366 
	,N9367,N9368,N9369,N9370,N9371,N9372,N9373,N9375 
	,N9376,N9377,N9378,N9379,N9380,N9381,N9383,N9384 
	,N9385,N9386,N9387,N9388,N9389,N9391,N9392,N9393 
	,N9394,N9396,N9397,N9398,N9399,N9400,N9401,N9402 
	,N9403,N9404,N9405,N9406,N9407,N9408,N9409,N9410 
	,N9411,N9413,N9414,N9415,N9416,N9417,N9418,N9419 
	,N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428 
	,N9430,N9431,N9432,N9433,N9434,N9435,N9436,N9437 
	,N9438,N9439,N9440,N9441,N9442,N9443,N9445,N9446 
	,N9447,N9448,N9449,N9450,N9451,N9453,N9454,N9455 
	,N9456,N9457,N9458,N9459,N9460,N9461,N9462,N9465 
	,N9466,N9467,N9468,N9469,N9470,N9471,N9472,N9473 
	,N9474,N9475,N9476,N9477,N9478,N9479,N9480,N9482 
	,N9483,N9484,N9485,N9486,N9487,N9490,N9491,N9492 
	,N9493,N9494,N9495,N9496,N9497,N9498,N9499,N9500 
	,N9501,N9502,N9503,N9504,N9505,N9507,N9508,N9509 
	,N9510,N9511,N9513,N9514,N9515,N9517,N9518,N9519 
	,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527 
	,N9528,N9529,N9530,N9531,N9532,N9533,N9534,N9535 
	,N9536,N9537,N9538,N9539,N9540,N9541,N9542,N9543 
	,N9545,N9546,N9547,N9548,N9549,N9551,N9552,N9553 
	,N9555,N9556,N9557,N9559,N9560,N9561,N9562,N9563 
	,N9564,N9565,N9566,N9567,N9568,N9569,N9570,N9571 
	,N9572,N9573,N9575,N9576,N9577,N9578,N9579,N9581 
	,N9582,N9583,N9585,N9586,N9587,N9588,N9589,N9590 
	,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598 
	,N9599,N9600,N9601,N9602,N9604,N9605,N9606,N9607 
	,N9608,N9609,N9610,N9611,N9612,N9613,N9614,N9615 
	,N9616,N9617,N9618,N9619,N9620,N9621,N9622,N9623 
	,N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632 
	,N9633,N9634,N9635,N9636,N9637,N9638,N9639,N9640 
	,N9642,N9643,N9644,N9645,N9646,N9647,N9648,N9650 
	,N9652,N9653,N9654,N9655,N9656,N9657,N9658,N9659 
	,N9660,N9661,N9662,N9663,N9664,N9665,N9666,N9667 
	,N9668,N9669,N9670,N9672,N9673,N9674,N9675,N9676 
	,N9677,N9678,N9680,N9681,N9682,N9683,N9684,N9685 
	,N9686,N9687,N9688,N9689,N9690,N9691,N9692,N9693 
	,N9694,N9695,N9696,N9697,N9698,N9699,N9700,N9701 
	,N9702,N9704,N9705,N9706,N9707,N9708,N9709,N9710 
	,N9712,N9714,N9715,N9716,N9717,N9718,N9719,N9720 
	,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728 
	,N9729,N9730,N9732,N9733,N9734,N9735,N9736,N9738 
	,N9739,N9741,N9742,N9743,N9744,N9745,N9746,N9747 
	,N9748,N9749,N9751,N9752,N9753,N9754,N9755,N9756 
	,N9757,N9759,N9760,N9761,N9762,N9763,N9764,N9765 
	,N9766,N9768,N9769,N9770,N9771,N9772,N9773,N9774 
	,N9775,N9776,N9778,N9779,N9780,N9781,N9782,N9784 
	,N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792 
	,N9793,N9794,N9796,N9797,N9798,N9799,N9800,N9801 
	,N9802,N9804,N9805,N9806,N9807,N9808,N9809,N9810 
	,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818 
	,N9819,N9821,N9822,N9823,N9824,N9825,N9826,N9827 
	,N9829,N9830,N9831,N9832,N9833,N9834,N9835,N9836 
	,N9837,N9838,N9839,N9840,N9841,N9842,N9843,N9845 
	,N9846,N9847,N9848,N9849,N9850,N9851,N9852,N9853 
	,N9854,N9855,N9856,N9857,N9859,N9860,N9861,N9862 
	,N9863,N9864,N9865,N9868,N9869,N9870,N9871,N9872 
	,N9873,N9874,N9875,N9876,N9877,N9878,N9879,N9880 
	,N9881,N9882,N9883,N9884,N9885,N9887,N9888,N9889 
	,N9890,N9891,N9893,N9894,N9895,N9896,N9897,N9898 
	,N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906 
	,N9907,N9908,N9909,N9910,N9911,N9912,N9913,N9914 
	,N9915,N9917,N9918,N9919,N9920,N9921,N9922,N9923 
	,N9924,N9925,N9927,N9928,N9929,N9930,N9932,N9933 
	,N9934,N9935,N9936,N9937,N9938,N9939,N9940,N9941 
	,N9942,N9944,N9945,N9946,N9947,N9949,N9950,N9952 
	,N9953,N9954,N9955,N9956,N9957,N9958,N9959,N9960 
	,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968 
	,N9969,N9970,N9971,N9973,N9974,N9975,N9976,N9977 
	,N9978,N9979,N9980,N9981,N9982,N9983,N9984,N9985 
	,N9986,N9987,N9988,N9989,N9990,N9991,N9993,N9994 
	,N9995,N9996,N9997,N9998,N9999,N10000,N10001,N10002 
	,N10003,N10004,N10005,N10007,N10008,N10009,N10010,N10011 
	,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021 
	,N10022,N10023,N10024,N10025,N10026,N10027,N10028,N10029 
	,N10030,N10031,N10032,N10033,N10034,N10035,N10037,N10038 
	,N10039,N10040,N10041,N10043,N10044,N10045,N10046,N10047 
	,N10048,N10049,N10050,N10051,N10052,N10053,N10054,N10055 
	,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10063 
	,N10064,N10066,N10067,N10068,N10071,N10072,N10073,N10074 
	,N10075,N10076,N10077,N10078,N10079,N10080,N10081,N10082 
	,N10083,N10084,N10085,N10086,N10087,N10088,N10089,N10090 
	,N10092,N10093,N10094,N10096,N10098,N10099,N10100,N10101 
	,N10102,N10103,N10104,N10105,N10106,N10107,N10108,N10110 
	,N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118 
	,N10119,N10120,N10121,N10122,N10123,N10124,N10125,N10126 
	,N10128,N10129,N10130,N10131,N10132,N10134,N10135,N10136 
	,N10137,N10138,N10140,N10141,N10142,N10143,N10144,N10145 
	,N10146,N10147,N10148,N10149,N10150,N10151,N10152,N10153 
	,N10155,N10156,N10157,N10158,N10160,N10161,N10163,N10164 
	,N10165,N10166,N10167,N10168,N10169,N10170,N10171,N10172 
	,N10173,N10174,N10175,N10176,N10177,N10178,N10179,N10180 
	,N10181,N10182,N10184,N10185,N10186,N10187,N10188,N10190 
	,N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198 
	,N10199,N10201,N10202,N10203,N10204,N10205,N10206,N10207 
	,N10208,N10209,N10210,N10211,N10212,N10214,N10215,N10216 
	,N10217,N10218,N10220,N10222,N10223,N10224,N10225,N10226 
	,N10227,N10228,N10229,N10230,N10231,N10232,N10233,N10234 
	,N10235,N10236,N10237,N10238,N10240,N11827,N11829,N11830 
	,N11833,N11834,N11836,N11837,N11838,N11839,N11840,N11843 
	,N11844,N11846,N11847,N11848,N11850,N11852,N11853,N11854 
	,N11856,N11858,N11859,N11863,N11864,N11865,N11866,N11867 
	,N11869,N11872,N11873,N11876,N11878,N11879,N11880,N11881 
	,N11885,N11886,N11887,N11888,N11889,N11890,N11892,N11893 
	,N11895,N11896,N11897,N11900,N11901,N11903,N11904,N11906 
	,N11909,N11910,N11911,N11912,N11913,N11915,N11916,N11919 
	,N11920,N11921,N11922,N11923,N11926,N11928,N11930,N11931 
	,N11933,N11934,N11935,N11937,N11941,N11942,N11943,N11944 
	,N11947,N11948,N11950,N11953,N11954,N11956,N11957,N11958 
	,N11960,N11963,N11964,N11965,N11966,N11967,N11969,N11971 
	,N11973,N11974,N11976,N11977,N11979,N11980,N11982,N11983 
	,N11985,N11986,N11987,N11988,N11990,N11992,N11993,N11995 
	,N11997,N11999,N12000,N12001,N12002,N12004,N12005,N12007 
	,N12010,N12011,N12012,N12014,N12016,N12019,N12021,N12023 
	,N12024,N12025,N12026,N12027,N12028,N12031,N12032,N12034 
	,N12035,N12037,N12038,N12040,N12041,N12042,N12044,N12045 
	,N12047,N12048,N12049,N12050,N12051,N12054,N12055,N12056 
	,N12057,N12059,N12061,N12062,N12063,N12065,N12066,N12068 
	,N12070,N12072,N12073,N12074,N12075,N12078,N12079,N12080 
	,N12081,N12082,N12083,N12084,N12086,N12087,N12089,N12090 
	,N12091,N12092,N12097,N12099,N12100,N12103,N12104,N12105 
	,N12106,N12108,N12111,N12112,N12114,N12115,N12116,N12117 
	,N12121,N12122,N12125,N12126,N12127,N12129,N12130,N12133 
	,N12134,N12136,N12137,N12138,N12141,N12142,N12144,N12145 
	,N12147,N12149,N12150,N12151,N12152,N12154,N12155,N12158 
	,N12159,N12160,N12161,N12162,N12165,N12166,N12168,N12169 
	,N12171,N12172,N12174,N12175,N12177,N12178,N12181,N12182 
	,N12183,N12184,N12187,N12188,N12190,N12191,N12193,N12194 
	,N12196,N12198,N12199,N12200,N12201,N12203,N12204,N12207 
	,N12208,N12210,N12212,N12213,N12215,N12216,N12218,N12219 
	,N12220,N12221,N12222,N12223,N12225,N12228,N12231,N12232 
	,N12234,N12235,N12238,N12239,N12241,N12242,N12243,N12244 
	,N12245,N12246,N12250,N12251,N12253,N12254,N12255,N12257 
	,N12259,N12261,N12262,N12265,N12267,N12268,N12269,N12270 
	,N12271,N12272,N12275,N12276,N12277,N12278,N12280,N12281 
	,N12283,N12285,N12287,N12288,N12291,N12293,N12294,N12295 
	,N12298,N12299,N12300,N12301,N12303,N12305,N12306,N12307 
	,N12309,N12310,N12311,N12314,N12316,N12317,N12318,N12321 
	,N12322,N12323,N12325,N12326,N12327,N12329,N12333,N12334 
	,N12335,N12336,N12340,N12341,N12343,N12344,N12345,N12347 
	,N12348,N12350,N12352,N12353,N12356,N12357,N12358,N12359 
	,N12360,N12363,N12364,N12365,N12367,N12368,N12370,N12372 
	,N12373,N12374,N12376,N12380,N12381,N12382,N12383,N12386 
	,N12387,N12388,N12390,N12391,N12393,N12394,N12396,N12399 
	,N12402,N12403,N12405,N12407,N12408,N12410,N12413,N12414 
	,N12416,N12417,N12418,N12419,N12422,N12425,N12426,N12427 
	,N12429,N12430,N12432,N12433,N12435,N12436,N12438,N12439 
	,N12440,N12442,N12443,N12444,N12445,N12448,N12449,N12452 
	,N13110,N13114,N13138,N13141,N13161,N13163,N13184,N13192 
	,N13195,N13197,N13201,N13203,N13206,N13212,N13216,N13270 
	,N13272,N13275,N13277,N13278,N13279,N13281,N13284,N13285 
	,N13286,N13287,N13289,N13290,N13292,N13293,N13294,N13296 
	,N13297,N13298,N13300,N13303,N13305,N13306,N13308,N13309 
	,N13311,N13312,N13313,N13314,N13315,N13317,N13318,N13321 
	,N13322,N13324,N13325,N13326,N13329,N13330,N13331,N13332 
	,N13333,N13335,N13336,N13337,N13340,N13342,N13343,N13344 
	,N13345,N13347,N13349,N13408,N13410,N13413,N13428,N13429 
	,N13430,N13433,N13434,N13435,N13436,N13439,N13440,N13441 
	,N13444,N13445,N13447,N13448,N13449,N13450,N13451,N13454 
	,N13455,N13456,N13459,N13460,N13463,N13464,N13465,N13466 
	,N13469,N13470,N13471,N13472,N13473,N13477,N13478,N13479 
	,N13480,N13483,N13484,N13485,N13486,N13487,N13489,N13491 
	,N13492,N13493,N13494,N13496,N13498,N13500,N13501,N13502 
	,N13503,N13504,N13507,N13508,N13509,N13512,N13513,N13514 
	,N13515,N13516,N13519,N13520,N13521,N13522,N13525,N13527 
	,N13529,N13532,N13533,N13534,N13535,N13536,N13539,N13540 
	,N13541,N13542,N13543,N13546,N13547,N13548,N13549,N13550 
	,N13553,N13554,N13555,N13556,N13559,N13560,N13561,N13565 
	,N13566,N13567,N13568,N13571,N13572,N13573,N13576,N13577 
	,N13578,N13757,N13872,N13897,N13910,N18828,N18830,N18832 
	,N18845,N18854,N18861,N18865,N18874,N37297;
INVXL inst_blk01_cellmath__39_I185 (.Y(N3966), .A(a_man[0]));
INVXL inst_blk01_cellmath__39_I186 (.Y(N4434), .A(a_man[1]));
INVXL inst_blk01_cellmath__39_I187 (.Y(N4398), .A(a_man[2]));
INVXL inst_blk01_cellmath__39_I188 (.Y(N4445), .A(a_man[3]));
INVXL inst_blk01_cellmath__39_I189 (.Y(N4304), .A(a_man[4]));
INVXL inst_blk01_cellmath__39_I190 (.Y(N4631), .A(a_man[5]));
INVXL inst_blk01_cellmath__39_I191 (.Y(N4097), .A(a_man[6]));
INVXL inst_blk01_cellmath__39_I192 (.Y(N4525), .A(a_man[7]));
INVXL inst_blk01_cellmath__39_I193 (.Y(N4121), .A(a_man[8]));
INVXL inst_blk01_cellmath__39_I194 (.Y(N4432), .A(a_man[9]));
INVXL inst_blk01_cellmath__39_I195 (.Y(N4032), .A(a_man[10]));
INVXL inst_blk01_cellmath__39_I196 (.Y(N4339), .A(a_man[11]));
INVXL inst_blk01_cellmath__39_I197 (.Y(N3939), .A(a_man[12]));
INVXL inst_blk01_cellmath__39_I198 (.Y(N4253), .A(a_man[13]));
INVXL inst_blk01_cellmath__39_I199 (.Y(N4565), .A(a_man[14]));
INVXL inst_blk01_cellmath__39_I200 (.Y(N4162), .A(a_man[15]));
INVXL inst_blk01_cellmath__39_I201 (.Y(N4471), .A(a_man[16]));
INVXL inst_blk01_cellmath__39_I202 (.Y(N4069), .A(a_man[17]));
INVXL inst_blk01_cellmath__39_I203 (.Y(N4385), .A(a_man[18]));
INVXL inst_blk01_cellmath__39_I204 (.Y(N3975), .A(a_man[19]));
INVXL inst_blk01_cellmath__39_I205 (.Y(N4291), .A(a_man[20]));
INVXL inst_blk01_cellmath__39_I206 (.Y(N4612), .A(a_man[21]));
INVXL inst_blk01_cellmath__39_I207 (.Y(N4198), .A(a_man[22]));
INVXL inst_blk01_cellmath__39_I208 (.Y(N4290), .A(N4445));
ADDHX1 inst_blk01_cellmath__39_I209 (.CO(N4352), .S(N4199), .A(N4304), .B(N4445));
ADDHX1 inst_blk01_cellmath__39_I210 (.CO(N3950), .S(N4513), .A(N4631), .B(N4398));
ADDFX1 inst_blk01_cellmath__39_I211 (.CO(N4174), .S(N4021), .A(N3966), .B(N4445), .CI(a_man[6]));
ADDHX1 inst_blk01_cellmath__39_I212 (.CO(N4484), .S(N4325), .A(N4525), .B(N4097));
ADDFX1 inst_blk01_cellmath__39_I213 (.CO(N4080), .S(N4652), .A(N4434), .B(N4304), .CI(N4325));
ADDHX1 inst_blk01_cellmath__39_I214 (.CO(N4396), .S(N4234), .A(N4121), .B(N4631));
ADDFX1 inst_blk01_cellmath__39_I215 (.CO(N3985), .S(N4548), .A(N4484), .B(N4398), .CI(N4234));
ADDFX1 inst_blk01_cellmath__39_I216 (.CO(N4456), .S(N4367), .A(N4097), .B(a_man[0]), .CI(N4432));
ADDFX1 inst_blk01_cellmath__39_I217 (.CO(N4301), .S(N4148), .A(N4445), .B(N4396), .CI(N4367));
ADDFX1 inst_blk01_cellmath__39_I218 (.CO(N4208), .S(N4250), .A(N4032), .B(a_man[1]), .CI(N4525));
ADDFX1 inst_blk01_cellmath__39_I219 (.CO(N4055), .S(N4628), .A(N4304), .B(N4456), .CI(N4250));
ADDFX1 inst_blk01_cellmath__39_I220 (.CO(N3962), .S(N4136), .A(N4121), .B(a_man[2]), .CI(N4339));
ADDFX1 inst_blk01_cellmath__39_I221 (.CO(N4522), .S(N4366), .A(N4631), .B(N4208), .CI(N4136));
ADDFX1 inst_blk01_cellmath__39_I222 (.CO(N4429), .S(N4015), .A(N3939), .B(a_man[3]), .CI(N4432));
ADDFX1 inst_blk01_cellmath__39_I223 (.CO(N4274), .S(N4117), .A(N3962), .B(N4097), .CI(N4015));
ADDFX1 inst_blk01_cellmath__39_I224 (.CO(N4184), .S(N4626), .A(N4253), .B(a_man[4]), .CI(N4032));
ADDFX1 inst_blk01_cellmath__39_I225 (.CO(N4030), .S(N4590), .A(N4525), .B(N4429), .CI(N4626));
XNOR2X1 inst_blk01_cellmath__39_I226 (.Y(N4337), .A(a_man[5]), .B(N3966));
OR2XL inst_blk01_cellmath__39_I227 (.Y(N4498), .A(a_man[5]), .B(N3966));
ADDFX1 inst_blk01_cellmath__39_I228 (.CO(N4560), .S(N3995), .A(N4339), .B(N4565), .CI(N4121));
ADDFX1 inst_blk01_cellmath__39_I229 (.CO(N4406), .S(N4248), .A(N4184), .B(N4337), .CI(N3995));
ADDFX1 inst_blk01_cellmath__39_I230 (.CO(N4160), .S(N3999), .A(N4434), .B(a_man[6]), .CI(N4162));
ADDFX1 inst_blk01_cellmath__39_I231 (.CO(N4639), .S(N4604), .A(N4432), .B(N3939), .CI(N4498));
ADDFX1 inst_blk01_cellmath__39_I232 (.CO(N4467), .S(N4313), .A(N4560), .B(N3999), .CI(N4604));
ADDHX1 inst_blk01_cellmath__39_I233 (.CO(N4219), .S(N4066), .A(a_man[7]), .B(N4398));
ADDFX1 inst_blk01_cellmath__39_I234 (.CO(N4536), .S(N4382), .A(N4471), .B(a_man[0]), .CI(N4253));
ADDFX1 inst_blk01_cellmath__39_I235 (.CO(N4287), .S(N4478), .A(N4066), .B(N4032), .CI(N4160));
ADDFX1 inst_blk01_cellmath__39_I236 (.CO(N4134), .S(N3972), .A(N4382), .B(N4639), .CI(N4478));
ADDFX1 inst_blk01_cellmath__39_I237 (.CO(N4041), .S(N4360), .A(N4445), .B(a_man[8]), .CI(N4069));
ADDFX1 inst_blk01_cellmath__39_I238 (.CO(N4608), .S(N4442), .A(N4219), .B(N4536), .CI(N4360));
ADDFX1 inst_blk01_cellmath__39_I239 (.CO(N4507), .S(N4242), .A(N4339), .B(a_man[1]), .CI(N4565));
ADDFX1 inst_blk01_cellmath__39_I240 (.CO(N4350), .S(N4194), .A(N4442), .B(N4287), .CI(N4242));
XNOR2X1 inst_blk01_cellmath__39_I241 (.Y(N3948), .A(a_man[9]), .B(N4304));
OR2XL inst_blk01_cellmath__39_I242 (.Y(N4104), .A(a_man[9]), .B(N4304));
ADDFX1 inst_blk01_cellmath__39_I243 (.CO(N4172), .S(N4343), .A(N4385), .B(a_man[2]), .CI(N4162));
ADDFX1 inst_blk01_cellmath__39_I244 (.CO(N4014), .S(N4573), .A(N4507), .B(N4041), .CI(N4343));
ADDFX1 inst_blk01_cellmath__39_I245 (.CO(N4649), .S(N4225), .A(N3966), .B(N3939), .CI(N3948));
ADDFX1 inst_blk01_cellmath__39_I246 (.CO(N4480), .S(N4322), .A(N4573), .B(N4608), .CI(N4225));
ADDFX1 inst_blk01_cellmath__39_I247 (.CO(N4230), .S(N4076), .A(N4631), .B(a_man[10]), .CI(N3975));
ADDFX1 inst_blk01_cellmath__39_I248 (.CO(N3984), .S(N4109), .A(N4471), .B(a_man[3]), .CI(N4253));
ADDFX1 inst_blk01_cellmath__39_I249 (.CO(N4546), .S(N4393), .A(N4172), .B(N4076), .CI(N4109));
ADDFX1 inst_blk01_cellmath__39_I250 (.CO(N4453), .S(N3988), .A(N4104), .B(N4434), .CI(N4649));
ADDFX1 inst_blk01_cellmath__39_I251 (.CO(N4298), .S(N4145), .A(N4014), .B(N4393), .CI(N3988));
ADDFX1 inst_blk01_cellmath__39_I252 (.CO(N4052), .S(N4624), .A(N4097), .B(a_man[11]), .CI(N4291));
ADDFX1 inst_blk01_cellmath__39_I253 (.CO(N4519), .S(N4592), .A(N4069), .B(a_man[4]), .CI(N4565));
ADDFX1 inst_blk01_cellmath__39_I254 (.CO(N4364), .S(N4206), .A(N3984), .B(N4624), .CI(N4592));
ADDFX1 inst_blk01_cellmath__39_I255 (.CO(N4271), .S(N4472), .A(N4230), .B(N4398), .CI(N4546));
ADDFX1 inst_blk01_cellmath__39_I256 (.CO(N4114), .S(N3958), .A(N4453), .B(N4206), .CI(N4472));
ADDFX1 inst_blk01_cellmath__39_I257 (.CO(N4586), .S(N4427), .A(N4525), .B(a_man[12]), .CI(N4612));
ADDFX1 inst_blk01_cellmath__39_I258 (.CO(N4335), .S(N4353), .A(N4162), .B(a_man[5]), .CI(N4385));
ADDFX1 inst_blk01_cellmath__39_I259 (.CO(N4182), .S(N4027), .A(N4519), .B(N4427), .CI(N4353));
ADDFX1 inst_blk01_cellmath__39_I260 (.CO(N4090), .S(N4235), .A(N4052), .B(N4445), .CI(N4364));
ADDFX1 inst_blk01_cellmath__39_I261 (.CO(N4658), .S(N4494), .A(N4027), .B(N4271), .CI(N4235));
ADDFX1 inst_blk01_cellmath__39_I262 (.CO(N4403), .S(N4244), .A(N4121), .B(a_man[13]), .CI(N4198));
ADDFX1 inst_blk01_cellmath__39_I263 (.CO(N4156), .S(N4116), .A(N3975), .B(a_man[6]), .CI(N4471));
ADDFX1 inst_blk01_cellmath__39_I264 (.CO(N3993), .S(N4556), .A(N4335), .B(N4116), .CI(N4244));
ADDFX1 inst_blk01_cellmath__39_I265 (.CO(N4636), .S(N4000), .A(N4586), .B(N4304), .CI(N4182));
ADDFX1 inst_blk01_cellmath__39_I266 (.CO(N4463), .S(N4309), .A(N4556), .B(N4090), .CI(N4000));
ADDFX1 inst_blk01_cellmath__39_I267 (.CO(N4214), .S(N4064), .A(N4291), .B(N4565), .CI(N4432));
ADDFX1 inst_blk01_cellmath__39_I268 (.CO(N4284), .S(N4574), .A(N4069), .B(a_man[7]), .CI(N4631));
ADDFX1 inst_blk01_cellmath__39_I269 (.CO(N4129), .S(N3969), .A(N4403), .B(N4156), .CI(N4574));
ADDFX1 inst_blk01_cellmath__39_I270 (.CO(N4037), .S(N4454), .A(N4064), .B(N3966), .CI(N3993));
ADDFX1 inst_blk01_cellmath__39_I271 (.CO(N4603), .S(N4438), .A(N4636), .B(N3969), .CI(N4454));
XNOR2X1 inst_blk01_cellmath__39_I272 (.Y(N4333), .A(a_man[15]), .B(N4032));
OR2XL inst_blk01_cellmath__39_I273 (.Y(N4505), .A(a_man[15]), .B(N4032));
ADDFX1 inst_blk01_cellmath__39_I274 (.CO(N4346), .S(N4191), .A(N4284), .B(N4214), .CI(N4333));
ADDFX1 inst_blk01_cellmath__39_I275 (.CO(N4258), .S(N4215), .A(N4612), .B(a_man[8]), .CI(N4385));
ADDFX1 inst_blk01_cellmath__39_I276 (.CO(N4100), .S(N3944), .A(N4434), .B(N4097), .CI(N4215));
ADDFX1 inst_blk01_cellmath__39_I277 (.CO(N4009), .S(N4101), .A(N4129), .B(a_man[14]), .CI(N4191));
ADDFX1 inst_blk01_cellmath__39_I278 (.CO(N4569), .S(N4414), .A(N3944), .B(N4037), .CI(N4101));
ADDFX1 inst_blk01_cellmath__39_I279 (.CO(N4320), .S(N4166), .A(N4198), .B(N4339), .CI(N4471));
ADDFX1 inst_blk01_cellmath__39_I280 (.CO(N4227), .S(N4073), .A(N3975), .B(a_man[9]), .CI(N4525));
ADDFX1 inst_blk01_cellmath__39_I281 (.CO(N3980), .S(N3953), .A(N4398), .B(a_man[0]), .CI(N4505));
ADDFX1 inst_blk01_cellmath__39_I282 (.CO(N4543), .S(N4388), .A(N4073), .B(N4166), .CI(N3953));
ADDFX1 inst_blk01_cellmath__39_I283 (.CO(N4449), .S(N4550), .A(N4346), .B(N4258), .CI(N4100));
ADDFX1 inst_blk01_cellmath__39_I284 (.CO(N4295), .S(N4141), .A(N4388), .B(N4009), .CI(N4550));
ADDFX1 inst_blk01_cellmath__39_I285 (.CO(N4049), .S(N4618), .A(N4291), .B(N3939), .CI(N4069));
ADDFX1 inst_blk01_cellmath__39_I286 (.CO(N3955), .S(N4516), .A(N4121), .B(a_man[10]), .CI(N4445));
ADDFX1 inst_blk01_cellmath__39_I287 (.CO(N4423), .S(N4410), .A(a_man[16]), .B(a_man[1]), .CI(N4227));
ADDFX1 inst_blk01_cellmath__39_I288 (.CO(N4268), .S(N4110), .A(N4618), .B(N3980), .CI(N4410));
ADDFX1 inst_blk01_cellmath__39_I289 (.CO(N4179), .S(N4293), .A(N4516), .B(N4320), .CI(N4543));
ADDFX1 inst_blk01_cellmath__39_I290 (.CO(N4024), .S(N4584), .A(N4449), .B(N4110), .CI(N4293));
ADDFX1 inst_blk01_cellmath__39_I291 (.CO(N4655), .S(N4175), .A(N4253), .B(a_man[18]), .CI(N4612));
ADDFX1 inst_blk01_cellmath__39_I292 (.CO(N4489), .S(N4331), .A(N3955), .B(N4049), .CI(N4175));
ADDFX1 inst_blk01_cellmath__39_I293 (.CO(N4400), .S(N4056), .A(N4304), .B(a_man[11]), .CI(N4432));
ADDFX1 inst_blk01_cellmath__39_I294 (.CO(N4238), .S(N4086), .A(a_man[17]), .B(a_man[2]), .CI(N4056));
ADDFX1 inst_blk01_cellmath__39_I295 (.CO(N4151), .S(N3937), .A(N4331), .B(N4423), .CI(N4086));
ADDFX1 inst_blk01_cellmath__39_I296 (.CO(N3989), .S(N4552), .A(N4268), .B(N4179), .CI(N3937));
ADDFX1 inst_blk01_cellmath__39_I297 (.CO(N4458), .S(N4306), .A(N4198), .B(N4565), .CI(N3975));
ADDFX1 inst_blk01_cellmath__39_I298 (.CO(N4372), .S(N4211), .A(N4032), .B(a_man[12]), .CI(N4631));
ADDFX1 inst_blk01_cellmath__39_I299 (.CO(N4124), .S(N4511), .A(a_man[0]), .B(a_man[3]), .CI(N4655));
ADDFX1 inst_blk01_cellmath__39_I300 (.CO(N3965), .S(N4527), .A(N4211), .B(N4306), .CI(N4511));
ADDFX1 inst_blk01_cellmath__39_I301 (.CO(N4597), .S(N4394), .A(N4489), .B(N4400), .CI(N4238));
ADDFX1 inst_blk01_cellmath__39_I302 (.CO(N4433), .S(N4280), .A(N4151), .B(N4527), .CI(N4394));
ADDFX1 inst_blk01_cellmath__39_I303 (.CO(N4187), .S(N4033), .A(N4339), .B(N4162), .CI(N4291));
ADDFX1 inst_blk01_cellmath__39_I304 (.CO(N4096), .S(N3940), .A(a_man[4]), .B(a_man[13]), .CI(N4097));
ADDFX1 inst_blk01_cellmath__39_I305 (.CO(N4566), .S(N4247), .A(a_man[19]), .B(a_man[1]), .CI(N4372));
ADDFX1 inst_blk01_cellmath__39_I306 (.CO(N4409), .S(N4255), .A(N4033), .B(N4124), .CI(N4247));
ADDFX1 inst_blk01_cellmath__39_I307 (.CO(N4317), .S(N4132), .A(N3940), .B(N4458), .CI(N3965));
ADDFX1 inst_blk01_cellmath__39_I308 (.CO(N4163), .S(N4005), .A(N4597), .B(N4255), .CI(N4132));
ADDHX1 inst_blk01_cellmath__39_I309 (.CO(N4641), .S(N4473), .A(a_man[21]), .B(N4471));
ADDFX1 inst_blk01_cellmath__39_I310 (.CO(N4386), .S(N4012), .A(N3939), .B(a_man[14]), .CI(N4525));
ADDFX1 inst_blk01_cellmath__39_I311 (.CO(N4224), .S(N4070), .A(N4096), .B(N4187), .CI(N4012));
ADDFX1 inst_blk01_cellmath__39_I312 (.CO(N4138), .S(N4621), .A(a_man[2]), .B(a_man[5]), .CI(a_man[0]));
ADDFX1 inst_blk01_cellmath__39_I313 (.CO(N3977), .S(N4541), .A(a_man[20]), .B(N4473), .CI(N4621));
ADDFX1 inst_blk01_cellmath__39_I314 (.CO(N4614), .S(N4493), .A(N4541), .B(N4566), .CI(N4070));
ADDFX1 inst_blk01_cellmath__39_I315 (.CO(N4447), .S(N4292), .A(N4409), .B(N4317), .CI(N4493));
XNOR2X1 inst_blk01_cellmath__39_I316 (.Y(N4046), .A(N4069), .B(N4253));
OR2XL inst_blk01_cellmath__39_I317 (.Y(N4200), .A(N4069), .B(N4253));
ADDFX1 inst_blk01_cellmath__39_I318 (.CO(N4266), .S(N4601), .A(a_man[15]), .B(a_man[22]), .CI(N4121));
ADDFX1 inst_blk01_cellmath__39_I319 (.CO(N4107), .S(N3952), .A(N4386), .B(N4046), .CI(N4601));
ADDFX1 inst_blk01_cellmath__39_I320 (.CO(N4023), .S(N4474), .A(a_man[3]), .B(a_man[6]), .CI(a_man[1]));
ADDFX1 inst_blk01_cellmath__39_I321 (.CO(N4581), .S(N4421), .A(N4641), .B(N4138), .CI(N4474));
ADDFX1 inst_blk01_cellmath__39_I322 (.CO(N4486), .S(N4355), .A(N4224), .B(N3977), .CI(N4421));
ADDFX1 inst_blk01_cellmath__39_I323 (.CO(N4326), .S(N4177), .A(N3952), .B(N4614), .CI(N4355));
ADDFX1 inst_blk01_cellmath__39_I324 (.CO(N4236), .S(N4237), .A(N4385), .B(a_man[16]), .CI(N4565));
ADDFX1 inst_blk01_cellmath__39_I325 (.CO(N4082), .S(N4653), .A(N4023), .B(N4266), .CI(N4237));
ADDFX1 inst_blk01_cellmath__39_I326 (.CO(N3987), .S(N4123), .A(N4432), .B(a_man[7]), .CI(a_man[4]));
ADDFX1 inst_blk01_cellmath__39_I327 (.CO(N4549), .S(N4397), .A(a_man[2]), .B(N4200), .CI(N4123));
ADDFX1 inst_blk01_cellmath__39_I328 (.CO(N4457), .S(N4004), .A(N4107), .B(N4581), .CI(N4653));
ADDFX1 inst_blk01_cellmath__39_I329 (.CO(N4302), .S(N4149), .A(N4397), .B(N4486), .CI(N4004));
ADDHX1 inst_blk01_cellmath__39_I330 (.CO(N4058), .S(N4630), .A(a_man[17]), .B(N3975));
ADDFX1 inst_blk01_cellmath__39_I331 (.CO(N4369), .S(N4210), .A(N4162), .B(a_man[8]), .CI(N4032));
ADDFX1 inst_blk01_cellmath__39_I332 (.CO(N4120), .S(N4613), .A(a_man[3]), .B(a_man[5]), .CI(N4630));
ADDFX1 inst_blk01_cellmath__39_I333 (.CO(N3963), .S(N4524), .A(N4236), .B(N4210), .CI(N4613));
ADDFX1 inst_blk01_cellmath__39_I334 (.CO(N4591), .S(N4485), .A(N4082), .B(N3987), .CI(N4549));
ADDFX1 inst_blk01_cellmath__39_I335 (.CO(N4430), .S(N4276), .A(N4457), .B(N4524), .CI(N4485));
ADDHX1 inst_blk01_cellmath__39_I336 (.CO(N4186), .S(N4031), .A(a_man[18]), .B(N4291));
ADDFX1 inst_blk01_cellmath__39_I337 (.CO(N4500), .S(N4338), .A(N4471), .B(a_man[9]), .CI(N4339));
ADDFX1 inst_blk01_cellmath__39_I338 (.CO(N4252), .S(N4368), .A(a_man[4]), .B(a_man[6]), .CI(N4058));
ADDFX1 inst_blk01_cellmath__39_I339 (.CO(N4093), .S(N3936), .A(N4338), .B(N4120), .CI(N4368));
ADDFX1 inst_blk01_cellmath__39_I340 (.CO(N4002), .S(N4249), .A(N4369), .B(N4031), .CI(N3963));
ADDFX1 inst_blk01_cellmath__39_I341 (.CO(N4562), .S(N4407), .A(N3936), .B(N4591), .CI(N4249));
ADDHX1 inst_blk01_cellmath__39_I342 (.CO(N4314), .S(N4161), .A(a_man[19]), .B(N4612));
ADDFX1 inst_blk01_cellmath__39_I343 (.CO(N4640), .S(N4470), .A(N4069), .B(a_man[10]), .CI(N3939));
ADDFX1 inst_blk01_cellmath__39_I344 (.CO(N4383), .S(N4135), .A(a_man[5]), .B(a_man[7]), .CI(N4186));
ADDFX1 inst_blk01_cellmath__39_I345 (.CO(N4221), .S(N4067), .A(N4470), .B(N4252), .CI(N4135));
ADDFX1 inst_blk01_cellmath__39_I346 (.CO(N4137), .S(N4016), .A(N4500), .B(N4161), .CI(N4093));
ADDFX1 inst_blk01_cellmath__39_I347 (.CO(N3974), .S(N4538), .A(N4067), .B(N4002), .CI(N4016));
ADDHX1 inst_blk01_cellmath__39_I348 (.CO(N4444), .S(N4288), .A(a_man[20]), .B(N4198));
ADDFX1 inst_blk01_cellmath__39_I349 (.CO(N4043), .S(N4609), .A(N4385), .B(a_man[11]), .CI(N4253));
ADDFX1 inst_blk01_cellmath__39_I350 (.CO(N4510), .S(N4625), .A(a_man[6]), .B(a_man[8]), .CI(N4314));
ADDFX1 inst_blk01_cellmath__39_I351 (.CO(N4351), .S(N4197), .A(N4609), .B(N4383), .CI(N4625));
ADDFX1 inst_blk01_cellmath__39_I352 (.CO(N4264), .S(N4495), .A(N4640), .B(N4288), .CI(N4221));
ADDFX1 inst_blk01_cellmath__39_I353 (.CO(N4105), .S(N3949), .A(N4197), .B(N4137), .CI(N4495));
ADDFX1 inst_blk01_cellmath__39_I354 (.CO(N4577), .S(N4420), .A(N3975), .B(a_man[21]), .CI(N4565));
ADDFX1 inst_blk01_cellmath__39_I355 (.CO(N4324), .S(N4377), .A(a_man[9]), .B(a_man[12]), .CI(a_man[7]));
ADDFX1 inst_blk01_cellmath__39_I356 (.CO(N4173), .S(N4018), .A(N4420), .B(N4510), .CI(N4377));
ADDFX1 inst_blk01_cellmath__39_I357 (.CO(N4078), .S(N4260), .A(N4043), .B(N4444), .CI(N4351));
ADDFX1 inst_blk01_cellmath__39_I358 (.CO(N4651), .S(N4482), .A(N4018), .B(N4264), .CI(N4260));
XNOR2X1 inst_blk01_cellmath__39_I359 (.Y(N4232), .A(N4291), .B(N4162));
OR2XL inst_blk01_cellmath__39_I360 (.Y(N4395), .A(N4291), .B(N4162));
ADDFX1 inst_blk01_cellmath__39_I361 (.CO(N4455), .S(N4359), .A(a_man[13]), .B(a_man[22]), .CI(a_man[10]));
ADDFX1 inst_blk01_cellmath__39_I362 (.CO(N4300), .S(N4147), .A(N4577), .B(N4232), .CI(N4359));
ADDFX1 inst_blk01_cellmath__39_I363 (.CO(N4207), .S(N4241), .A(N4324), .B(a_man[8]), .CI(N4173));
ADDFX1 inst_blk01_cellmath__39_I364 (.CO(N4053), .S(N4627), .A(N4147), .B(N4078), .CI(N4241));
ADDFX1 inst_blk01_cellmath__39_I365 (.CO(N3960), .S(N4126), .A(N4612), .B(a_man[14]), .CI(N4471));
ADDFX1 inst_blk01_cellmath__39_I366 (.CO(N4521), .S(N4365), .A(N4395), .B(N4455), .CI(N4126));
ADDFX1 inst_blk01_cellmath__39_I367 (.CO(N4428), .S(N4006), .A(a_man[9]), .B(a_man[11]), .CI(N4300));
ADDFX1 inst_blk01_cellmath__39_I368 (.CO(N4273), .S(N4115), .A(N4365), .B(N4207), .CI(N4006));
ADDHX1 inst_blk01_cellmath__39_I369 (.CO(N4029), .S(N4588), .A(a_man[15]), .B(N4198));
ADDFX1 inst_blk01_cellmath__39_I370 (.CO(N4336), .S(N4183), .A(a_man[10]), .B(a_man[12]), .CI(N4069));
ADDFX1 inst_blk01_cellmath__39_I371 (.CO(N4092), .S(N4617), .A(N3960), .B(N4588), .CI(N4183));
ADDFX1 inst_blk01_cellmath__39_I372 (.CO(N3934), .S(N4496), .A(N4428), .B(N4521), .CI(N4617));
ADDFX1 inst_blk01_cellmath__39_I373 (.CO(N4404), .S(N4246), .A(N4385), .B(a_man[16]), .CI(a_man[13]));
ADDFX1 inst_blk01_cellmath__39_I374 (.CO(N4158), .S(N4488), .A(N4336), .B(a_man[11]), .CI(N4029));
ADDFX1 inst_blk01_cellmath__39_I375 (.CO(N3996), .S(N4557), .A(N4246), .B(N4092), .CI(N4488));
XNOR2X1 inst_blk01_cellmath__39_I376 (.Y(N4311), .A(N3975), .B(a_man[17]));
OR2XL inst_blk01_cellmath__39_I377 (.Y(N4466), .A(N3975), .B(a_man[17]));
ADDFX1 inst_blk01_cellmath__39_I378 (.CO(N4533), .S(N4594), .A(a_man[12]), .B(a_man[14]), .CI(N4404));
ADDFX1 inst_blk01_cellmath__39_I379 (.CO(N4378), .S(N4218), .A(N4311), .B(N4158), .CI(N4594));
XNOR2X1 inst_blk01_cellmath__39_I380 (.Y(N3970), .A(N4291), .B(a_man[18]));
OR2XL inst_blk01_cellmath__39_I381 (.Y(N4130), .A(N4291), .B(a_man[18]));
ADDFX1 inst_blk01_cellmath__39_I382 (.CO(N4193), .S(N3976), .A(a_man[13]), .B(a_man[15]), .CI(N4466));
ADDFX1 inst_blk01_cellmath__39_I383 (.CO(N4039), .S(N4605), .A(N3970), .B(N4533), .CI(N3976));
XNOR2X1 inst_blk01_cellmath__39_I384 (.Y(N4348), .A(N4612), .B(a_man[19]));
OR2XL inst_blk01_cellmath__39_I385 (.Y(N4506), .A(N4612), .B(a_man[19]));
ADDFX1 inst_blk01_cellmath__39_I386 (.CO(N4571), .S(N4081), .A(a_man[14]), .B(a_man[16]), .CI(N4130));
ADDFX1 inst_blk01_cellmath__39_I387 (.CO(N4417), .S(N4262), .A(N4348), .B(N4193), .CI(N4081));
XNOR2X1 inst_blk01_cellmath__39_I388 (.Y(N4011), .A(N4198), .B(a_man[20]));
OR2XL inst_blk01_cellmath__39_I389 (.Y(N4170), .A(N4198), .B(a_man[20]));
ADDFX1 inst_blk01_cellmath__39_I390 (.CO(N4229), .S(N4185), .A(a_man[15]), .B(a_man[17]), .CI(N4506));
ADDFX1 inst_blk01_cellmath__39_I391 (.CO(N4075), .S(N4647), .A(N4011), .B(N4571), .CI(N4185));
ADDFX1 inst_blk01_cellmath__39_I392 (.CO(N4545), .S(N4391), .A(a_man[16]), .B(a_man[18]), .CI(N4612));
ADDFX1 inst_blk01_cellmath__39_I393 (.CO(N4451), .S(N4297), .A(N4229), .B(N4170), .CI(N4391));
ADDFX1 inst_blk01_cellmath__39_I394 (.CO(N4204), .S(N4042), .A(a_man[19]), .B(a_man[22]), .CI(a_man[17]));
ADDFX1 inst_blk01_cellmath__39_I395 (.CO(N4051), .S(N4622), .A(a_man[21]), .B(N4545), .CI(N4042));
ADDFX1 inst_blk01_cellmath__39_I396 (.CO(N4518), .S(N4361), .A(a_man[18]), .B(a_man[20]), .CI(N4204));
ADDHX1 inst_blk01_cellmath__39_I397 (.CO(N4112), .S(N3957), .A(a_man[21]), .B(a_man[19]));
ADDHX1 inst_blk01_cellmath__39_I398 (.CO(N4425), .S(N4270), .A(a_man[22]), .B(a_man[20]));
INVXL inst_blk01_cellmath__39_I399 (.Y(N4088), .A(N4398));
NOR2XL inst_blk01_cellmath__39_I400 (.Y(N4243), .A(N3966), .B(N4290));
NAND2XL inst_blk01_cellmath__39_I401 (.Y(N4402), .A(N3966), .B(N4290));
NOR2XL inst_blk01_cellmath__39_I402 (.Y(N4554), .A(N4434), .B(N4199));
NAND2XL inst_blk01_cellmath__39_I403 (.Y(N3992), .A(N4434), .B(N4199));
NOR2XL inst_blk01_cellmath__39_I404 (.Y(N4154), .A(N4513), .B(N4352));
NAND2XL inst_blk01_cellmath__39_I405 (.Y(N4308), .A(N4352), .B(N4513));
AND2XL inst_blk01_cellmath__39_I407 (.Y(N4634), .A(N3950), .B(N4021));
NOR2XL inst_blk01_cellmath__39_I408 (.Y(N4062), .A(N4174), .B(N4652));
NAND2XL inst_blk01_cellmath__39_I409 (.Y(N4213), .A(N4174), .B(N4652));
AND2XL inst_blk01_cellmath__39_I411 (.Y(N4530), .A(N4080), .B(N4548));
NOR2XL inst_blk01_cellmath__39_I412 (.Y(N3968), .A(N3985), .B(N4148));
NAND2XL inst_blk01_cellmath__39_I413 (.Y(N4127), .A(N3985), .B(N4148));
NOR2XL inst_blk01_cellmath__39_I414 (.Y(N4282), .A(N4301), .B(N4628));
NAND2XL inst_blk01_cellmath__39_I415 (.Y(N4437), .A(N4301), .B(N4628));
NOR2XL inst_blk01_cellmath__39_I416 (.Y(N4599), .A(N4055), .B(N4366));
NOR2XL inst_blk01_cellmath__39_I418 (.Y(N4190), .A(N4522), .B(N4117));
NAND2XL inst_blk01_cellmath__39_I419 (.Y(N4344), .A(N4522), .B(N4117));
NOR2XL inst_blk01_cellmath__39_I420 (.Y(N4503), .A(N4274), .B(N4590));
NOR2XL inst_blk01_cellmath__39_I422 (.Y(N4098), .A(N4030), .B(N4248));
NAND2XL inst_blk01_cellmath__39_I423 (.Y(N4256), .A(N4030), .B(N4248));
NOR2XL inst_blk01_cellmath__39_I424 (.Y(N4413), .A(N4406), .B(N4313));
NAND2XL inst_blk01_cellmath__39_I425 (.Y(N4567), .A(N4406), .B(N4313));
NOR2XL inst_blk01_cellmath__39_I426 (.Y(N4007), .A(N4467), .B(N3972));
NAND2XL inst_blk01_cellmath__39_I427 (.Y(N4165), .A(N4467), .B(N3972));
NOR2XL inst_blk01_cellmath__39_I428 (.Y(N4318), .A(N4134), .B(N4194));
NOR2XL inst_blk01_cellmath__39_I430 (.Y(N4643), .A(N4350), .B(N4322));
NAND2XL inst_blk01_cellmath__39_I431 (.Y(N4071), .A(N4350), .B(N4322));
NOR2XL inst_blk01_cellmath__39_I432 (.Y(N3978), .A(a_man[1]), .B(a_man[0]));
AOI21XL inst_blk01_cellmath__39_I433 (.Y(N4047), .A0(N4402), .A1(N4088), .B0(N4243));
INVXL inst_blk01_cellmath__39_I434 (.Y(N4201), .A(N4402));
OAI21XL inst_blk01_cellmath__39_I435 (.Y(N4329), .A0(N4201), .A1(N3978), .B0(N4047));
AO21XL inst_blk01_cellmath__39_I436 (.Y(N4514), .A0(N4308), .A1(N4554), .B0(N4154));
AOI31X1 inst_blk01_cellmath__39_I438 (.Y(N4595), .A0(N4308), .A1(N3992), .A2(N4329), .B0(N4514));
OAI22XL inst_blk01_cellmath__39_I8318 (.Y(N4222), .A0(N4634), .A1(N4595), .B0(N3950), .B1(N4021));
AOI21XL inst_blk01_cellmath__39_I442 (.Y(N4580), .A0(N4213), .A1(N4222), .B0(N4062));
OAI22XL inst_blk01_cellmath__39_I8319 (.Y(N4118), .A0(N4530), .A1(N4580), .B0(N4080), .B1(N4548));
AO21XL inst_blk01_cellmath__39_I446 (.Y(N4563), .A0(N4437), .A1(N3968), .B0(N4282));
AOI31X1 inst_blk01_cellmath__39_I448 (.Y(N4508), .A0(N4437), .A1(N4127), .A2(N4118), .B0(N4563));
AOI21XL inst_blk01_cellmath__39_I449 (.Y(N4418), .A0(N4344), .A1(N4599), .B0(N4190));
OAI2BB1X1 inst_blk01_cellmath__39_I8320 (.Y(N4576), .A0N(N4055), .A1N(N4366), .B0(N4344));
AOI21XL inst_blk01_cellmath__39_I452 (.Y(N4323), .A0(N4256), .A1(N4503), .B0(N4098));
OAI2BB1X1 inst_blk01_cellmath__39_I8321 (.Y(N4481), .A0N(N4274), .A1N(N4590), .B0(N4256));
OAI21XL inst_blk01_cellmath__39_I457 (.Y(N4600), .A0(N4481), .A1(N4418), .B0(N4323));
NOR3XL inst_blk01_cellmath__39_I458 (.Y(N4283), .A(N4481), .B(N4576), .C(N4508));
OR2XL inst_blk01_cellmath__39_I459 (.Y(N4347), .A(N4283), .B(N4600));
AO21XL inst_blk01_cellmath__39_I460 (.Y(N3961), .A0(N4165), .A1(N4413), .B0(N4007));
AOI31X1 inst_blk01_cellmath__39_I467 (.Y(N4460), .A0(N4165), .A1(N4567), .A2(N4347), .B0(N3961));
AOI21XL inst_blk01_cellmath__39_I470 (.Y(N4373), .A0(N4071), .A1(N4318), .B0(N4643));
OAI2BB1X1 inst_blk01_cellmath__39_I8322 (.Y(N4529), .A0N(N4134), .A1N(N4194), .B0(N4071));
OAI21XL inst_blk01_cellmath__39_I473 (.Y(N3935), .A0(N4529), .A1(N4460), .B0(N4373));
NOR2XL inst_blk01_cellmath__39_I509 (.Y(N4559), .A(N4298), .B(N3958));
XOR2XL inst_blk01_cellmath__39_I510 (.Y(N4001), .A(N4298), .B(N3958));
XOR2XL inst_blk01_cellmath__39_I511 (.Y(N4312), .A(N4114), .B(N4494));
NOR2XL inst_blk01_cellmath__39_I512 (.Y(N4468), .A(N4658), .B(N4309));
XOR2XL inst_blk01_cellmath__39_I513 (.Y(N4638), .A(N4658), .B(N4309));
XOR2XL inst_blk01_cellmath__39_I514 (.Y(N4220), .A(N4463), .B(N4438));
NOR2XL inst_blk01_cellmath__39_I515 (.Y(N4381), .A(N4603), .B(N4414));
XOR2XL inst_blk01_cellmath__39_I516 (.Y(N4535), .A(N4603), .B(N4414));
XOR2XL inst_blk01_cellmath__39_I517 (.Y(N4133), .A(N4569), .B(N4141));
NOR2XL inst_blk01_cellmath__39_I518 (.Y(N4286), .A(N4295), .B(N4584));
XOR2XL inst_blk01_cellmath__39_I519 (.Y(N4443), .A(N4295), .B(N4584));
XOR2XL inst_blk01_cellmath__39_I520 (.Y(N4040), .A(N4024), .B(N4552));
NOR2XL inst_blk01_cellmath__39_I521 (.Y(N4195), .A(N3989), .B(N4280));
XOR2XL inst_blk01_cellmath__39_I522 (.Y(N4349), .A(N3989), .B(N4280));
XOR2XL inst_blk01_cellmath__39_I523 (.Y(N3947), .A(N4433), .B(N4005));
NOR2XL inst_blk01_cellmath__39_I524 (.Y(N4103), .A(N4163), .B(N4292));
XOR2XL inst_blk01_cellmath__39_I525 (.Y(N4263), .A(N4163), .B(N4292));
XOR2XL inst_blk01_cellmath__39_I526 (.Y(N4575), .A(N4447), .B(N4177));
NOR2XL inst_blk01_cellmath__39_I527 (.Y(N4013), .A(N4326), .B(N4149));
XOR2XL inst_blk01_cellmath__39_I528 (.Y(N4171), .A(N4326), .B(N4149));
XOR2XL inst_blk01_cellmath__39_I529 (.Y(N4479), .A(N4302), .B(N4276));
NOR2XL inst_blk01_cellmath__39_I530 (.Y(N4648), .A(N4430), .B(N4407));
XOR2XL inst_blk01_cellmath__39_I531 (.Y(N4077), .A(N4430), .B(N4407));
XOR2XL inst_blk01_cellmath__39_I532 (.Y(N4392), .A(N4562), .B(N4538));
NOR2XL inst_blk01_cellmath__39_I533 (.Y(N4547), .A(N3974), .B(N3949));
XOR2XL inst_blk01_cellmath__39_I534 (.Y(N3983), .A(N3974), .B(N3949));
XOR2XL inst_blk01_cellmath__39_I535 (.Y(N4299), .A(N4105), .B(N4482));
NOR2XL inst_blk01_cellmath__39_I536 (.Y(N4452), .A(N4651), .B(N4627));
XOR2XL inst_blk01_cellmath__39_I537 (.Y(N4623), .A(N4651), .B(N4627));
XOR2XL inst_blk01_cellmath__39_I538 (.Y(N4205), .A(N4053), .B(N4115));
NOR2XL inst_blk01_cellmath__39_I539 (.Y(N4363), .A(N4273), .B(N4496));
XOR2XL inst_blk01_cellmath__39_I540 (.Y(N4520), .A(N4273), .B(N4496));
XOR2XL inst_blk01_cellmath__39_I541 (.Y(N4113), .A(N4557), .B(N3934));
NOR2XL inst_blk01_cellmath__39_I542 (.Y(N4272), .A(N3996), .B(N4218));
XOR2XL inst_blk01_cellmath__39_I543 (.Y(N4426), .A(N3996), .B(N4218));
XOR2XL inst_blk01_cellmath__39_I544 (.Y(N4028), .A(N4378), .B(N4605));
NOR2XL inst_blk01_cellmath__39_I545 (.Y(N4181), .A(N4039), .B(N4262));
XOR2XL inst_blk01_cellmath__39_I546 (.Y(N4334), .A(N4039), .B(N4262));
XOR2XL inst_blk01_cellmath__39_I547 (.Y(N4657), .A(N4417), .B(N4647));
NOR2XL inst_blk01_cellmath__39_I548 (.Y(N4089), .A(N4297), .B(N4075));
XOR2XL inst_blk01_cellmath__39_I549 (.Y(N4245), .A(N4297), .B(N4075));
XOR2XL inst_blk01_cellmath__39_I550 (.Y(N4555), .A(N4451), .B(N4622));
NOR2XL inst_blk01_cellmath__39_I551 (.Y(N3994), .A(N4361), .B(N4051));
XOR2XL inst_blk01_cellmath__39_I552 (.Y(N4155), .A(N4361), .B(N4051));
XOR2XL inst_blk01_cellmath__39_I553 (.Y(N4464), .A(N3957), .B(N4518));
NOR2XL inst_blk01_cellmath__39_I554 (.Y(N4635), .A(N4112), .B(N4270));
XOR2XL inst_blk01_cellmath__39_I555 (.Y(N4063), .A(N4112), .B(N4270));
XOR2XL inst_blk01_cellmath__39_I556 (.Y(N4376), .A(N4612), .B(N4425));
XNOR2X1 inst_blk01_cellmath__39_I557 (.Y(N4169), .A(a_man[22]), .B(a_man[21]));
INVXL cmpii_A_I8384 (.Y(N18830), .A(N4480));
INVXL cmpii_A_I8385 (.Y(N18832), .A(N4145));
AND2XL cmpii_A_I8386 (.Y(N18828), .A(N18830), .B(N18832));
OAI22XL cmpii_A_I8387 (.Y(N4128), .A0(N18828), .A1(N3935), .B0(N18830), .B1(N18832));
AOI2BB2X1 inst_blk01_cellmath__39_I559 (.Y(N4439), .A0N(N4114), .A1N(N4494), .B0(N4559), .B1(N4312));
NAND2XL inst_blk01_cellmath__39_I560 (.Y(N4602), .A(N4312), .B(N4001));
AOI2BB2X1 inst_blk01_cellmath__39_I561 (.Y(N4036), .A0N(N4463), .A1N(N4438), .B0(N4468), .B1(N4220));
NAND2XL inst_blk01_cellmath__39_I562 (.Y(N4192), .A(N4220), .B(N4638));
AOI2BB2X1 inst_blk01_cellmath__39_I563 (.Y(N4345), .A0N(N4569), .A1N(N4141), .B0(N4381), .B1(N4133));
NAND2XL inst_blk01_cellmath__39_I564 (.Y(N4504), .A(N4133), .B(N4535));
AOI2BB2X1 inst_blk01_cellmath__39_I565 (.Y(N3945), .A0N(N4024), .A1N(N4552), .B0(N4286), .B1(N4040));
NAND2XL inst_blk01_cellmath__39_I566 (.Y(N4099), .A(N4040), .B(N4443));
AOI2BB2X1 inst_blk01_cellmath__39_I567 (.Y(N4257), .A0N(N4433), .A1N(N4005), .B0(N4195), .B1(N3947));
NAND2XL inst_blk01_cellmath__39_I568 (.Y(N4415), .A(N3947), .B(N4349));
AOI2BB2X1 inst_blk01_cellmath__39_I569 (.Y(N4568), .A0N(N4447), .A1N(N4177), .B0(N4103), .B1(N4575));
NAND2XL inst_blk01_cellmath__39_I570 (.Y(N4008), .A(N4575), .B(N4263));
AOI2BB2X1 inst_blk01_cellmath__39_I571 (.Y(N4167), .A0N(N4302), .A1N(N4276), .B0(N4013), .B1(N4479));
NAND2XL inst_blk01_cellmath__39_I572 (.Y(N4319), .A(N4479), .B(N4171));
AOI2BB2X1 inst_blk01_cellmath__39_I573 (.Y(N4476), .A0N(N4562), .A1N(N4538), .B0(N4648), .B1(N4392));
NAND2XL inst_blk01_cellmath__39_I574 (.Y(N4645), .A(N4392), .B(N4077));
AOI2BB2X1 inst_blk01_cellmath__39_I575 (.Y(N4072), .A0N(N4105), .A1N(N4482), .B0(N4547), .B1(N4299));
NAND2XL inst_blk01_cellmath__39_I576 (.Y(N4226), .A(N4299), .B(N3983));
AOI2BB2X1 inst_blk01_cellmath__39_I577 (.Y(N4389), .A0N(N4053), .A1N(N4115), .B0(N4452), .B1(N4205));
NAND2XL inst_blk01_cellmath__39_I578 (.Y(N4542), .A(N4205), .B(N4623));
AOI2BB2X1 inst_blk01_cellmath__39_I579 (.Y(N3979), .A0N(N4557), .A1N(N3934), .B0(N4363), .B1(N4113));
NAND2XL inst_blk01_cellmath__39_I580 (.Y(N4142), .A(N4113), .B(N4520));
AOI2BB2X1 inst_blk01_cellmath__39_I581 (.Y(N4294), .A0N(N4378), .A1N(N4605), .B0(N4272), .B1(N4028));
NAND2XL inst_blk01_cellmath__39_I582 (.Y(N4448), .A(N4028), .B(N4426));
AOI2BB2X1 inst_blk01_cellmath__39_I583 (.Y(N4619), .A0N(N4417), .A1N(N4647), .B0(N4181), .B1(N4657));
NAND2XL inst_blk01_cellmath__39_I584 (.Y(N4048), .A(N4657), .B(N4334));
AOI2BB2X1 inst_blk01_cellmath__39_I585 (.Y(N4202), .A0N(N4451), .A1N(N4622), .B0(N4089), .B1(N4555));
NAND2XL inst_blk01_cellmath__39_I586 (.Y(N4356), .A(N4555), .B(N4245));
AOI2BB2X1 inst_blk01_cellmath__39_I587 (.Y(N4515), .A0N(N3957), .A1N(N4518), .B0(N3994), .B1(N4464));
NAND2XL inst_blk01_cellmath__39_I588 (.Y(N3954), .A(N4464), .B(N4155));
OAI21XL inst_blk01_cellmath__39_I589 (.Y(N4422), .A0(N4602), .A1(N4128), .B0(N4439));
OAI21XL inst_blk01_cellmath__39_I590 (.Y(N4025), .A0(N4504), .A1(N4036), .B0(N4345));
NOR2XL inst_blk01_cellmath__39_I591 (.Y(N4178), .A(N4504), .B(N4192));
OAI21XL inst_blk01_cellmath__39_I592 (.Y(N4330), .A0(N4415), .A1(N3945), .B0(N4257));
NOR2XL inst_blk01_cellmath__39_I593 (.Y(N4490), .A(N4415), .B(N4099));
OAI21XL inst_blk01_cellmath__39_I594 (.Y(N4654), .A0(N4319), .A1(N4568), .B0(N4167));
NOR2XL inst_blk01_cellmath__39_I595 (.Y(N4085), .A(N4319), .B(N4008));
OAI21XL inst_blk01_cellmath__39_I596 (.Y(N4239), .A0(N4226), .A1(N4476), .B0(N4072));
NOR2XL inst_blk01_cellmath__39_I597 (.Y(N4399), .A(N4226), .B(N4645));
OAI21XL inst_blk01_cellmath__39_I598 (.Y(N4551), .A0(N4142), .A1(N4389), .B0(N3979));
NOR2XL inst_blk01_cellmath__39_I599 (.Y(N3990), .A(N4142), .B(N4542));
OAI21XL inst_blk01_cellmath__39_I600 (.Y(N4150), .A0(N4048), .A1(N4294), .B0(N4619));
NOR2XL inst_blk01_cellmath__39_I601 (.Y(N4305), .A(N4048), .B(N4448));
OAI21XL inst_blk01_cellmath__39_I602 (.Y(N4459), .A0(N3954), .A1(N4202), .B0(N4515));
NOR2XL inst_blk01_cellmath__39_I603 (.Y(N4632), .A(N3954), .B(N4356));
AOI21XL inst_blk01_cellmath__39_I604 (.Y(N4059), .A0(N4178), .A1(N4422), .B0(N4025));
AOI21XL inst_blk01_cellmath__39_I605 (.Y(N4371), .A0(N4085), .A1(N4330), .B0(N4654));
NAND2XL inst_blk01_cellmath__39_I606 (.Y(N4526), .A(N4085), .B(N4490));
AOI21XL inst_blk01_cellmath__39_I607 (.Y(N4279), .A0(N4632), .A1(N4150), .B0(N4459));
NAND2XL inst_blk01_cellmath__39_I608 (.Y(N4435), .A(N4632), .B(N4305));
OAI21XL inst_blk01_cellmath__39_I609 (.Y(N4596), .A0(N4526), .A1(N4059), .B0(N4371));
AO21XL inst_blk01_cellmath__39_I610 (.Y(N4341), .A0(N3990), .A1(N4239), .B0(N4551));
AOI31X1 inst_blk01_cellmath__39_I611 (.Y(N4501), .A0(N3990), .A1(N4399), .A2(N4596), .B0(N4341));
INVXL inst_blk01_cellmath__39_I612 (.Y(N4095), .A(N4490));
INVXL inst_blk01_cellmath__39_I613 (.Y(N4254), .A(N4330));
OAI21XL inst_blk01_cellmath__39_I614 (.Y(N4411), .A0(N4095), .A1(N4059), .B0(N4254));
INVXL inst_blk01_cellmath__39_I615 (.Y(N4065), .A(N4596));
AOI21XL inst_blk01_cellmath__39_I616 (.Y(N4316), .A0(N4399), .A1(N4596), .B0(N4239));
INVXL inst_blk01_cellmath__39_I617 (.Y(N4216), .A(N4501));
INVXL inst_blk01_cellmath__39_I618 (.Y(N4223), .A(N4305));
INVXL inst_blk01_cellmath__39_I619 (.Y(N4387), .A(N4150));
OAI21XL inst_blk01_cellmath__39_I620 (.Y(N4540), .A0(N4223), .A1(N4501), .B0(N4387));
OAI21XL inst_blk01_cellmath__39_I621 (.Y(N4139), .A0(N4435), .A1(N4501), .B0(N4279));
INVXL inst_blk01_cellmath__39_I622 (.Y(N4446), .A(N4192));
INVXL inst_blk01_cellmath__39_I623 (.Y(N4615), .A(N4036));
AOI21XL inst_blk01_cellmath__39_I624 (.Y(N4045), .A0(N4446), .A1(N4422), .B0(N4615));
INVXL inst_blk01_cellmath__39_I625 (.Y(N4379), .A(N4059));
OAI21XL inst_blk01_cellmath__39_I626 (.Y(N3951), .A0(N4099), .A1(N4059), .B0(N3945));
INVXL inst_blk01_cellmath__39_I627 (.Y(N4534), .A(N4411));
INVXL inst_blk01_cellmath__39_I628 (.Y(N4582), .A(N4008));
INVXL inst_blk01_cellmath__39_I629 (.Y(N4022), .A(N4568));
AOI21XL inst_blk01_cellmath__39_I630 (.Y(N4176), .A0(N4582), .A1(N4411), .B0(N4022));
INVXL inst_blk01_cellmath__39_I631 (.Y(N3971), .A(N4065));
OAI21XL inst_blk01_cellmath__39_I632 (.Y(N4083), .A0(N4645), .A1(N4065), .B0(N4476));
INVXL inst_blk01_cellmath__39_I633 (.Y(N4131), .A(N4316));
OAI21XL inst_blk01_cellmath__39_I634 (.Y(N3986), .A0(N4542), .A1(N4316), .B0(N4389));
INVXL inst_blk01_cellmath__39_I635 (.Y(N4285), .A(N4216));
INVXL inst_blk01_cellmath__39_I636 (.Y(N4629), .A(N4448));
INVXL inst_blk01_cellmath__39_I637 (.Y(N4057), .A(N4294));
AOI21XL inst_blk01_cellmath__39_I638 (.Y(N4209), .A0(N4629), .A1(N4216), .B0(N4057));
INVXL inst_blk01_cellmath__39_I639 (.Y(N4441), .A(N4540));
INVXL inst_blk01_cellmath__39_I640 (.Y(N4119), .A(N4356));
INVXL inst_blk01_cellmath__39_I641 (.Y(N4275), .A(N4202));
AOI21XL inst_blk01_cellmath__39_I642 (.Y(N4431), .A0(N4119), .A1(N4540), .B0(N4275));
INVXL inst_blk01_cellmath__39_I643 (.Y(N4606), .A(N4139));
OAI2BB2XL inst_blk01_cellmath__39_I644 (.Y(N4499), .A0N(N4635), .A1N(N4376), .B0(N4612), .B1(N4425));
AOI31X1 inst_blk01_cellmath__39_I645 (.Y(N3938), .A0(N4376), .A1(N4063), .A2(N4139), .B0(N4499));
INVXL inst_blk01_cellmath__39_I650 (.Y(N4384), .A(N4535));
INVXL inst_blk01_cellmath__39_I651 (.Y(N4537), .A(N4381));
OAI21XL inst_blk01_cellmath__39_I652 (.Y(N3973), .A0(N4384), .A1(N4045), .B0(N4537));
AOI21XL inst_blk01_cellmath__39_I653 (.Y(N4611), .A0(N4443), .A1(N4379), .B0(N4286));
AOI21XL inst_blk01_cellmath__39_I654 (.Y(N4509), .A0(N4349), .A1(N3951), .B0(N4195));
INVXL inst_blk01_cellmath__39_I655 (.Y(N4419), .A(N4263));
INVXL inst_blk01_cellmath__39_I656 (.Y(N4579), .A(N4103));
OAI21XL inst_blk01_cellmath__39_I657 (.Y(N4017), .A0(N4419), .A1(N4534), .B0(N4579));
INVXL inst_blk01_cellmath__39_I658 (.Y(N4650), .A(N4171));
INVXL inst_blk01_cellmath__39_I659 (.Y(N4079), .A(N4013));
OAI21XL inst_blk01_cellmath__39_I660 (.Y(N4231), .A0(N4650), .A1(N4176), .B0(N4079));
AOI21XL inst_blk01_cellmath__39_I661 (.Y(N4146), .A0(N4077), .A1(N3971), .B0(N4648));
AOI21XL inst_blk01_cellmath__39_I662 (.Y(N4054), .A0(N3983), .A1(N4083), .B0(N4547));
AOI21XL inst_blk01_cellmath__39_I663 (.Y(N3959), .A0(N4623), .A1(N4131), .B0(N4452));
AOI21XL inst_blk01_cellmath__39_I664 (.Y(N4587), .A0(N4520), .A1(N3986), .B0(N4363));
INVXL inst_blk01_cellmath__39_I665 (.Y(N4497), .A(N4426));
INVXL inst_blk01_cellmath__39_I666 (.Y(N3933), .A(N4272));
OAI21XL inst_blk01_cellmath__39_I667 (.Y(N4091), .A0(N4497), .A1(N4285), .B0(N3933));
INVXL inst_blk01_cellmath__39_I668 (.Y(N3998), .A(N4334));
INVXL inst_blk01_cellmath__39_I669 (.Y(N4157), .A(N4181));
OAI21XL inst_blk01_cellmath__39_I670 (.Y(N4310), .A0(N3998), .A1(N4209), .B0(N4157));
INVXL inst_blk01_cellmath__39_I671 (.Y(N4217), .A(N4245));
INVXL inst_blk01_cellmath__39_I672 (.Y(N4380), .A(N4089));
OAI21XL inst_blk01_cellmath__39_I673 (.Y(N4532), .A0(N4217), .A1(N4441), .B0(N4380));
INVXL inst_blk01_cellmath__39_I674 (.Y(N4440), .A(N4155));
INVXL inst_blk01_cellmath__39_I675 (.Y(N4607), .A(N3994));
OAI21XL inst_blk01_cellmath__39_I676 (.Y(N4038), .A0(N4440), .A1(N4431), .B0(N4607));
INVXL inst_blk01_cellmath__39_I677 (.Y(N3946), .A(N4063));
INVXL inst_blk01_cellmath__39_I678 (.Y(N4102), .A(N4635));
OAI21XL inst_blk01_cellmath__39_I679 (.Y(N4261), .A0(N3946), .A1(N4606), .B0(N4102));
XNOR2X1 inst_blk01_cellmath__39_I686 (.Y(N623), .A(N3973), .B(N4133));
XNOR2X1 inst_blk01_cellmath__39_I687 (.Y(N624), .A(N4379), .B(N4443));
XOR2XL inst_blk01_cellmath__39_I688 (.Y(N625), .A(N4611), .B(N4040));
XNOR2X1 inst_blk01_cellmath__39_I689 (.Y(N626), .A(N3951), .B(N4349));
XOR2XL inst_blk01_cellmath__39_I690 (.Y(N627), .A(N4509), .B(N3947));
XOR2XL inst_blk01_cellmath__39_I691 (.Y(N628), .A(N4534), .B(N4263));
XNOR2X1 inst_blk01_cellmath__39_I692 (.Y(N629), .A(N4017), .B(N4575));
XOR2XL inst_blk01_cellmath__39_I693 (.Y(N630), .A(N4176), .B(N4171));
XNOR2X1 inst_blk01_cellmath__39_I694 (.Y(N631), .A(N4231), .B(N4479));
XNOR2X1 inst_blk01_cellmath__39_I695 (.Y(N632), .A(N3971), .B(N4077));
XOR2XL inst_blk01_cellmath__39_I696 (.Y(N633), .A(N4146), .B(N4392));
XNOR2X1 inst_blk01_cellmath__39_I697 (.Y(N634), .A(N4083), .B(N3983));
XOR2XL inst_blk01_cellmath__39_I698 (.Y(N635), .A(N4054), .B(N4299));
XNOR2X1 inst_blk01_cellmath__39_I699 (.Y(N636), .A(N4131), .B(N4623));
XOR2XL inst_blk01_cellmath__39_I700 (.Y(N637), .A(N3959), .B(N4205));
XNOR2X1 inst_blk01_cellmath__39_I701 (.Y(N638), .A(N3986), .B(N4520));
XOR2XL inst_blk01_cellmath__39_I702 (.Y(N639), .A(N4587), .B(N4113));
XOR2XL inst_blk01_cellmath__39_I703 (.Y(N640), .A(N4285), .B(N4426));
XNOR2X1 inst_blk01_cellmath__39_I704 (.Y(N641), .A(N4091), .B(N4028));
XOR2XL inst_blk01_cellmath__39_I705 (.Y(N642), .A(N4209), .B(N4334));
XNOR2X1 inst_blk01_cellmath__39_I706 (.Y(N643), .A(N4310), .B(N4657));
XOR2XL inst_blk01_cellmath__39_I707 (.Y(N644), .A(N4441), .B(N4245));
XNOR2X1 inst_blk01_cellmath__39_I708 (.Y(N645), .A(N4532), .B(N4555));
XOR2XL inst_blk01_cellmath__39_I709 (.Y(N646), .A(N4431), .B(N4155));
XNOR2X1 inst_blk01_cellmath__39_I710 (.Y(N647), .A(N4038), .B(N4464));
XOR2XL inst_blk01_cellmath__39_I711 (.Y(N648), .A(N4606), .B(N4063));
XNOR2X1 inst_blk01_cellmath__39_I712 (.Y(N649), .A(N4261), .B(N4376));
XNOR2X1 inst_blk01_cellmath__39_I713 (.Y(N650), .A(N3938), .B(N4169));
OA22X1 inst_blk01_cellmath__39_I714 (.Y(N652), .A0(N4169), .A1(N3938), .B0(a_man[22]), .B1(a_man[21]));
INVXL inst_blk01_cellmath__39_I715 (.Y(N651), .A(N652));
INVXL inst_cellmath__42_0_I717 (.Y(N5364), .A(a_exp[1]));
INVXL inst_cellmath__42_0_I718 (.Y(N5385), .A(a_exp[3]));
NAND2BXL inst_cellmath__42_0_I719 (.Y(N5373), .AN(N5364), .B(a_exp[2]));
NAND2XL inst_cellmath__42_0_I720 (.Y(N5372), .A(N5385), .B(N5373));
OR2XL inst_cellmath__42_0_I721 (.Y(N5371), .A(a_exp[4]), .B(N5372));
OR2XL inst_cellmath__42_0_I722 (.Y(N5379), .A(a_exp[5]), .B(N5371));
NOR2XL inst_cellmath__42_0_I723 (.Y(N5376), .A(a_exp[6]), .B(N5379));
INVXL inst_cellmath__42_0_I724 (.Y(inst_cellmath__42[1]), .A(N5364));
XOR2XL inst_cellmath__42_0_I727 (.Y(inst_cellmath__42[4]), .A(N5372), .B(a_exp[4]));
XOR2XL inst_cellmath__42_0_I729 (.Y(inst_cellmath__42[6]), .A(N5379), .B(a_exp[6]));
XOR2XL inst_cellmath__42_0_I730 (.Y(inst_cellmath__42[7]), .A(N5376), .B(a_exp[7]));
NOR2BX1 inst_cellmath__42_0_I731 (.Y(inst_cellmath__42[8]), .AN(a_exp[7]), .B(N5376));
MXI2XL inst_cellmath__48_I733 (.Y(N5438), .A(N624), .B(N623), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I734 (.Y(N5486), .A(N625), .B(N624), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I735 (.Y(N5534), .A(N626), .B(N625), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I736 (.Y(N5581), .A(N627), .B(N626), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I737 (.Y(N5411), .A(N628), .B(N627), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I738 (.Y(N5459), .A(N629), .B(N628), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I739 (.Y(N5507), .A(N630), .B(N629), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I740 (.Y(N5553), .A(N631), .B(N630), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I741 (.Y(N5601), .A(N632), .B(N631), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I742 (.Y(N5431), .A(N633), .B(N632), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I743 (.Y(N5479), .A(N634), .B(N633), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I744 (.Y(N5527), .A(N635), .B(N634), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I745 (.Y(N5574), .A(N636), .B(N635), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I746 (.Y(N5405), .A(N637), .B(N636), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I747 (.Y(N5450), .A(N638), .B(N637), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I748 (.Y(N5499), .A(N639), .B(N638), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I749 (.Y(N5546), .A(N640), .B(N639), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I750 (.Y(N5594), .A(N641), .B(N640), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I751 (.Y(N5425), .A(N642), .B(N641), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I752 (.Y(N5473), .A(N643), .B(N642), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I753 (.Y(N5519), .A(N644), .B(N643), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I754 (.Y(N5565), .A(N645), .B(N644), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I755 (.Y(N5612), .A(N646), .B(N645), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I756 (.Y(N5443), .A(N647), .B(N646), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I757 (.Y(N5491), .A(N648), .B(N647), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I758 (.Y(N5540), .A(N649), .B(N648), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I759 (.Y(N5585), .A(N650), .B(N649), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I760 (.Y(N5416), .A(N651), .B(N650), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I761 (.Y(N5464), .A(N652), .B(N651), .S0(a_exp[0]));
NAND2XL inst_cellmath__48_I762 (.Y(N5512), .A(N652), .B(a_exp[0]));
INVXL buf1_A_I23544 (.Y(N37297), .A(inst_cellmath__42[1]));
INVXL buf1_A_I23545 (.Y(N5451), .A(N37297));
MXI2XL inst_cellmath__48_I764 (.Y(N5478), .A(N5438), .B(N5534), .S0(N5451));
MXI2XL inst_cellmath__48_I765 (.Y(N5526), .A(N5486), .B(N5581), .S0(N5451));
MXI2XL inst_cellmath__48_I766 (.Y(N5571), .A(N5534), .B(N5411), .S0(N5451));
MXI2XL inst_cellmath__48_I767 (.Y(N5403), .A(N5581), .B(N5459), .S0(N5451));
MXI2XL inst_cellmath__48_I768 (.Y(N5449), .A(N5411), .B(N5507), .S0(N5451));
MXI2XL inst_cellmath__48_I769 (.Y(N5498), .A(N5459), .B(N5553), .S0(N5451));
MXI2XL inst_cellmath__48_I770 (.Y(N5545), .A(N5507), .B(N5601), .S0(N5451));
MXI2XL inst_cellmath__48_I771 (.Y(N5592), .A(N5553), .B(N5431), .S0(N5451));
MXI2XL inst_cellmath__48_I772 (.Y(N5422), .A(N5601), .B(N5479), .S0(N5451));
MXI2XL inst_cellmath__48_I773 (.Y(N5471), .A(N5431), .B(N5527), .S0(N5451));
MXI2XL inst_cellmath__48_I774 (.Y(N5518), .A(N5479), .B(N5574), .S0(N5451));
MXI2XL inst_cellmath__48_I775 (.Y(N5564), .A(N5527), .B(N5405), .S0(N5451));
MXI2XL inst_cellmath__48_I776 (.Y(N5611), .A(N5574), .B(N5450), .S0(N5451));
MXI2XL inst_cellmath__48_I777 (.Y(N5442), .A(N5405), .B(N5499), .S0(N5451));
MXI2XL inst_cellmath__48_I778 (.Y(N5489), .A(N5450), .B(N5546), .S0(N5451));
MXI2XL inst_cellmath__48_I779 (.Y(N5538), .A(N5499), .B(N5594), .S0(N5451));
MXI2XL inst_cellmath__48_I780 (.Y(N5584), .A(N5546), .B(N5425), .S0(N5451));
MXI2XL inst_cellmath__48_I781 (.Y(N5415), .A(N5594), .B(N5473), .S0(N5451));
MXI2XL inst_cellmath__48_I782 (.Y(N5462), .A(N5425), .B(N5519), .S0(N5451));
MXI2XL inst_cellmath__48_I783 (.Y(N5511), .A(N5473), .B(N5565), .S0(N5451));
MXI2XL inst_cellmath__48_I784 (.Y(N5557), .A(N5519), .B(N5612), .S0(N5451));
MXI2XL inst_cellmath__48_I785 (.Y(N5605), .A(N5565), .B(N5443), .S0(N5451));
MXI2XL inst_cellmath__48_I786 (.Y(N5434), .A(N5612), .B(N5491), .S0(N5451));
MXI2XL inst_cellmath__48_I787 (.Y(N5482), .A(N5443), .B(N5540), .S0(N5451));
MXI2XL inst_cellmath__48_I788 (.Y(N5531), .A(N5491), .B(N5585), .S0(N5451));
MXI2XL inst_cellmath__48_I789 (.Y(N5577), .A(N5540), .B(N5416), .S0(N5451));
MXI2XL inst_cellmath__48_I790 (.Y(N5409), .A(N5585), .B(N5464), .S0(N5451));
MXI2XL inst_cellmath__48_I791 (.Y(N5455), .A(N5416), .B(N5512), .S0(N5451));
NOR2XL inst_cellmath__48_I792 (.Y(N5504), .A(N5464), .B(N5451));
NOR2XL inst_cellmath__48_I793 (.Y(N5598), .A(N5512), .B(N5451));
CLKXOR2X1 inst_cellmath__48_I8324 (.Y(N5500), .A(inst_cellmath__42[1]), .B(a_exp[2]));
MXI2XL inst_cellmath__48_I795 (.Y(N5562), .A(N5449), .B(N5478), .S0(N5500));
MXI2XL inst_cellmath__48_I796 (.Y(N5610), .A(N5498), .B(N5526), .S0(N5500));
MXI2XL inst_cellmath__48_I797 (.Y(N5441), .A(N5545), .B(N5571), .S0(N5500));
MXI2XL inst_cellmath__48_I798 (.Y(N5487), .A(N5592), .B(N5403), .S0(N5500));
MXI2XL inst_cellmath__48_I799 (.Y(N5535), .A(N5422), .B(N5449), .S0(N5500));
MXI2XL inst_cellmath__48_I800 (.Y(N5583), .A(N5471), .B(N5498), .S0(N5500));
MXI2XL inst_cellmath__48_I801 (.Y(N5413), .A(N5518), .B(N5545), .S0(N5500));
MXI2XL inst_cellmath__48_I802 (.Y(N5461), .A(N5564), .B(N5592), .S0(N5500));
MXI2XL inst_cellmath__48_I803 (.Y(N5510), .A(N5611), .B(N5422), .S0(N5500));
MXI2XL inst_cellmath__48_I804 (.Y(N5554), .A(N5442), .B(N5471), .S0(N5500));
MXI2XL inst_cellmath__48_I805 (.Y(N5602), .A(N5489), .B(N5518), .S0(N5500));
MXI2XL inst_cellmath__48_I806 (.Y(N5433), .A(N5538), .B(N5564), .S0(N5500));
MXI2XL inst_cellmath__48_I807 (.Y(N5481), .A(N5584), .B(N5611), .S0(N5500));
MXI2XL inst_cellmath__48_I808 (.Y(N5530), .A(N5415), .B(N5442), .S0(N5500));
MXI2XL inst_cellmath__48_I809 (.Y(N5576), .A(N5462), .B(N5489), .S0(N5500));
MXI2XL inst_cellmath__48_I810 (.Y(N5406), .A(N5511), .B(N5538), .S0(N5500));
MXI2XL inst_cellmath__48_I811 (.Y(N5453), .A(N5557), .B(N5584), .S0(N5500));
MXI2XL inst_cellmath__48_I812 (.Y(N5503), .A(N5605), .B(N5415), .S0(N5500));
MXI2XL inst_cellmath__48_I813 (.Y(N5549), .A(N5434), .B(N5462), .S0(N5500));
MXI2XL inst_cellmath__48_I814 (.Y(N5597), .A(N5482), .B(N5511), .S0(N5500));
MXI2XL inst_cellmath__48_I815 (.Y(N5427), .A(N5531), .B(N5557), .S0(N5500));
MXI2XL inst_cellmath__48_I816 (.Y(N5474), .A(N5577), .B(N5605), .S0(N5500));
MXI2XL inst_cellmath__48_I817 (.Y(N5521), .A(N5409), .B(N5434), .S0(N5500));
MXI2XL inst_cellmath__48_I818 (.Y(N5568), .A(N5455), .B(N5482), .S0(N5500));
MXI2XL inst_cellmath__48_I819 (.Y(N5615), .A(N5504), .B(N5531), .S0(N5500));
MXI2XL inst_cellmath__48_I820 (.Y(N5446), .A(N5598), .B(N5577), .S0(N5500));
NAND2XL inst_cellmath__48_I821 (.Y(N5493), .A(N5409), .B(N5500));
NAND2XL inst_cellmath__48_I822 (.Y(N5587), .A(N5455), .B(N5500));
NAND2XL inst_cellmath__48_I823 (.Y(N5467), .A(N5504), .B(N5500));
NAND2XL inst_cellmath__48_I824 (.Y(N5560), .A(N5598), .B(N5500));
CLKXOR2X1 inst_cellmath__48_I8325 (.Y(N5593), .A(N5373), .B(N5385));
MXI2XL inst_cellmath__48_I826 (.Y(N5528), .A(N5562), .B(N5510), .S0(N5593));
MXI2XL inst_cellmath__48_I827 (.Y(N5573), .A(N5610), .B(N5554), .S0(N5593));
MXI2XL inst_cellmath__48_I828 (.Y(N5404), .A(N5441), .B(N5602), .S0(N5593));
MXI2XL inst_cellmath__48_I829 (.Y(N5452), .A(N5487), .B(N5433), .S0(N5593));
MXI2XL inst_cellmath__48_I830 (.Y(N5501), .A(N5535), .B(N5481), .S0(N5593));
MXI2XL inst_cellmath__48_I831 (.Y(N5547), .A(N5583), .B(N5530), .S0(N5593));
MXI2XL inst_cellmath__48_I832 (.Y(N5595), .A(N5413), .B(N5576), .S0(N5593));
MXI2XL inst_cellmath__48_I833 (.Y(N5424), .A(N5461), .B(N5406), .S0(N5593));
MXI2XL inst_cellmath__48_I834 (.Y(N5472), .A(N5510), .B(N5453), .S0(N5593));
MXI2XL inst_cellmath__48_I835 (.Y(N5520), .A(N5554), .B(N5503), .S0(N5593));
MXI2XL inst_cellmath__48_I836 (.Y(N5566), .A(N5602), .B(N5549), .S0(N5593));
MXI2XL inst_cellmath__48_I837 (.Y(N5613), .A(N5433), .B(N5597), .S0(N5593));
MXI2XL inst_cellmath__48_I838 (.Y(N5444), .A(N5481), .B(N5427), .S0(N5593));
MXI2XL inst_cellmath__48_I839 (.Y(N5490), .A(N5530), .B(N5474), .S0(N5593));
MXI2XL inst_cellmath__48_I840 (.Y(N5539), .A(N5576), .B(N5521), .S0(N5593));
MXI2XL inst_cellmath__48_I841 (.Y(N5586), .A(N5406), .B(N5568), .S0(N5593));
MXI2XL inst_cellmath__48_I842 (.Y(N5417), .A(N5453), .B(N5615), .S0(N5593));
MXI2XL inst_cellmath__48_I843 (.Y(N5465), .A(N5503), .B(N5446), .S0(N5593));
MXI2XL inst_cellmath__48_I844 (.Y(N5513), .A(N5549), .B(N5493), .S0(N5593));
MXI2XL inst_cellmath__48_I845 (.Y(N5558), .A(N5597), .B(N5587), .S0(N5593));
MXI2XL inst_cellmath__48_I846 (.Y(N5606), .A(N5427), .B(N5467), .S0(N5593));
MXI2XL inst_cellmath__48_I847 (.Y(N5436), .A(N5474), .B(N5560), .S0(N5593));
NOR2XL inst_cellmath__48_I848 (.Y(N5483), .A(N5521), .B(N5593));
NOR2XL inst_cellmath__48_I849 (.Y(N5578), .A(N5568), .B(N5593));
NOR2XL inst_cellmath__48_I850 (.Y(N5456), .A(N5615), .B(N5593));
NOR2XL inst_cellmath__48_I851 (.Y(N5550), .A(N5446), .B(N5593));
NOR2XL inst_cellmath__48_I852 (.Y(N5428), .A(N5493), .B(N5593));
NOR2XL inst_cellmath__48_I853 (.Y(N5523), .A(N5587), .B(N5593));
NOR2XL inst_cellmath__48_I854 (.Y(N5616), .A(N5467), .B(N5593));
NOR2XL inst_cellmath__48_I855 (.Y(N5494), .A(N5560), .B(N5593));
XNOR2X1 inst_cellmath__48_I8326 (.Y(N5423), .A(N5371), .B(a_exp[5]));
NAND2XL inst_cellmath__48_I857 (.Y(N5463), .A(N5528), .B(N5423));
NAND2XL inst_cellmath__48_I858 (.Y(N5556), .A(N5573), .B(N5423));
NAND2XL inst_cellmath__48_I859 (.Y(N5435), .A(N5404), .B(N5423));
NAND2XL inst_cellmath__48_I860 (.Y(N5532), .A(N5452), .B(N5423));
NAND2XL inst_cellmath__48_I861 (.Y(N5408), .A(N5501), .B(N5423));
NAND2XL inst_cellmath__48_I862 (.Y(N5505), .A(N5547), .B(N5423));
NAND2XL inst_cellmath__48_I863 (.Y(N5599), .A(N5595), .B(N5423));
NAND2XL inst_cellmath__48_I864 (.Y(N5476), .A(N5424), .B(N5423));
NAND2XL inst_cellmath__48_I865 (.Y(N5569), .A(N5472), .B(N5423));
NAND2XL inst_cellmath__48_I866 (.Y(N5447), .A(N5520), .B(N5423));
NAND2XL inst_cellmath__48_I867 (.Y(N5542), .A(N5566), .B(N5423));
NAND2XL inst_cellmath__48_I868 (.Y(N5419), .A(N5613), .B(N5423));
NAND2XL inst_cellmath__48_I869 (.Y(N5515), .A(N5444), .B(N5423));
NAND2XL inst_cellmath__48_I870 (.Y(N5608), .A(N5490), .B(N5423));
NAND2XL inst_cellmath__48_I871 (.Y(N5485), .A(N5539), .B(N5423));
NAND2XL inst_cellmath__48_I872 (.Y(N5580), .A(N5586), .B(N5423));
NAND2XL inst_cellmath__48_I873 (.Y(N5458), .A(N5417), .B(N5423));
NAND2XL inst_cellmath__48_I874 (.Y(N5552), .A(N5465), .B(N5423));
NAND2XL inst_cellmath__48_I875 (.Y(N5430), .A(N5513), .B(N5423));
NAND2XL inst_cellmath__48_I876 (.Y(N5525), .A(N5558), .B(N5423));
NAND2XL inst_cellmath__48_I877 (.Y(N5402), .A(N5606), .B(N5423));
NAND2XL inst_cellmath__48_I878 (.Y(N5497), .A(N5436), .B(N5423));
NAND2XL inst_cellmath__48_I879 (.Y(N5591), .A(N5483), .B(N5423));
NAND2XL inst_cellmath__48_I880 (.Y(N5470), .A(N5578), .B(N5423));
NAND2XL inst_cellmath__48_I881 (.Y(N5563), .A(N5456), .B(N5423));
NAND2XL inst_cellmath__48_I882 (.Y(N5440), .A(N5550), .B(N5423));
NAND2XL inst_cellmath__48_I883 (.Y(N5537), .A(N5428), .B(N5423));
NAND2XL inst_cellmath__48_I884 (.Y(N5414), .A(N5523), .B(N5423));
NAND2XL inst_cellmath__48_I885 (.Y(N5509), .A(N5616), .B(N5423));
NAND2XL inst_cellmath__48_I886 (.Y(N5604), .A(N5494), .B(N5423));
MXI2XL inst_cellmath__48_I887 (.Y(N684), .A(N5463), .B(N5458), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I888 (.Y(N685), .A(N5556), .B(N5552), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I889 (.Y(N686), .A(N5435), .B(N5430), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I890 (.Y(N687), .A(N5532), .B(N5525), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I891 (.Y(N688), .A(N5408), .B(N5402), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I892 (.Y(N689), .A(N5505), .B(N5497), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I893 (.Y(N690), .A(N5599), .B(N5591), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I894 (.Y(N691), .A(N5476), .B(N5470), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I895 (.Y(N692), .A(N5569), .B(N5563), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I896 (.Y(N693), .A(N5447), .B(N5440), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I897 (.Y(N694), .A(N5542), .B(N5537), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I898 (.Y(N695), .A(N5419), .B(N5414), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I899 (.Y(N696), .A(N5515), .B(N5509), .S0(inst_cellmath__42[4]));
MXI2XL inst_cellmath__48_I900 (.Y(N697), .A(N5608), .B(N5604), .S0(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I901 (.Y(N698), .A(N5485), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I902 (.Y(N699), .A(N5580), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I903 (.Y(N700), .A(N5458), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I904 (.Y(N701), .A(N5552), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I905 (.Y(N702), .A(N5430), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I906 (.Y(N703), .A(N5525), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I907 (.Y(N704), .A(N5402), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I908 (.Y(N705), .A(N5497), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I909 (.Y(N706), .A(N5591), .B(inst_cellmath__42[4]));
OR2XL inst_cellmath__48_I910 (.Y(N707), .A(N5470), .B(inst_cellmath__42[4]));
NOR2XL inst_cellmath__48_I911 (.Y(N708), .A(N5563), .B(inst_cellmath__42[4]));
XNOR2X1 cynw_cm_float_cos_I913 (.Y(N493), .A(N708), .B(N707));
INVXL inst_cellmath__61_0_I914 (.Y(N5817), .A(N707));
XNOR2X1 inst_cellmath__61_0_I916 (.Y(inst_cellmath__61[1]), .A(N685), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I917 (.Y(inst_cellmath__61[2]), .A(N686), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I918 (.Y(inst_cellmath__61[3]), .A(N687), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I919 (.Y(inst_cellmath__61[4]), .A(N688), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I920 (.Y(inst_cellmath__61[5]), .A(N689), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I921 (.Y(inst_cellmath__61[6]), .A(N690), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I922 (.Y(inst_cellmath__61[7]), .A(N691), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I923 (.Y(inst_cellmath__61[8]), .A(N692), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I924 (.Y(inst_cellmath__61[9]), .A(N693), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I925 (.Y(inst_cellmath__61[10]), .A(N694), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I926 (.Y(inst_cellmath__61[11]), .A(N695), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I927 (.Y(inst_cellmath__61[12]), .A(N696), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I928 (.Y(inst_cellmath__61[13]), .A(N697), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I929 (.Y(inst_cellmath__61[14]), .A(N698), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I930 (.Y(inst_cellmath__61[15]), .A(N699), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I932 (.Y(inst_cellmath__61[17]), .A(N701), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I933 (.Y(inst_cellmath__61[18]), .A(N702), .B(N5817));
XNOR2X1 inst_cellmath__61_0_I937 (.Y(inst_cellmath__61[22]), .A(N706), .B(N5817));
XOR2XL cynw_cm_float_cos_I8327 (.Y(inst_cellmath__115__W1[0]), .A(N700), .B(N5817));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I938 (.Y(N6011), .A(inst_cellmath__61[17]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I939 (.Y(N6139), .A(inst_cellmath__61[18]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I940 (.Y(N5877), .A(inst_cellmath__61[18]), .B(N6011));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I941 (.Y(N6198), .A(N6139), .B(N6011));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I942 (.Y(N6501), .A(N6139), .B(N6011));
AOI22X1 inst_cellmath__195__80__2WWMM_2WWMM_I943 (.Y(N6490), .A0(inst_cellmath__61[17]), .A1(inst_cellmath__61[18]), .B0(N6139), .B1(N6011));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I944 (.Y(N6411), .A(inst_cellmath__61[18]), .B(inst_cellmath__61[17]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I945 (.Y(N6021), .A(N6139), .B(inst_cellmath__61[17]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I946 (.Y(N6328), .A(N6139), .B(inst_cellmath__61[17]));
AOI22X1 inst_cellmath__195__80__2WWMM_2WWMM_I947 (.Y(N6241), .A0(N6011), .A1(inst_cellmath__61[18]), .B0(N6139), .B1(inst_cellmath__61[17]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I948 (.Y(N6238), .A(inst_cellmath__61[17]), .B(inst_cellmath__61[18]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I949 (.Y(N6487), .A(N6011), .B(inst_cellmath__61[18]));
XNOR2X4 inst_cellmath__195__80__2WWMM_2WWMM_I8328 (.Y(N6349), .A(N703), .B(N5817));
INVX3 inst_cellmath__195__80__2WWMM_2WWMM_I952 (.Y(N6273), .A(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I953 (.Y(N5928), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I954 (.Y(N6094), .A0(N6273), .A1(N6328), .B0(N5877), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I955 (.Y(N6147), .A(N6273), .B(N6139));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I956 (.Y(N5996), .A0(N6273), .A1(N6328), .B0(inst_cellmath__61[17]), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I957 (.Y(N6154), .A(N6273), .B(N6021));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I958 (.Y(N6448), .A0(N6273), .A1(N6490), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I959 (.Y(N5898), .A0(N6273), .A1(N6241), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I960 (.Y(N6059), .A0(N6273), .A1(N6021), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I961 (.Y(N6218), .A0(N6273), .A1(N6011), .B0(N6501), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I962 (.Y(N6370), .A(N6273), .B(N6328));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I963 (.Y(N5966), .A0(N6273), .A1(N5877), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I964 (.Y(N6365), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(inst_cellmath__61[18]), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I965 (.Y(N6281), .A(N6349), .B(N6139));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I966 (.Y(N5959), .A(N6273), .B(N6139));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I967 (.Y(N6343), .A0(N6273), .A1(N6490), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I968 (.Y(N6492), .A0(N6273), .A1(N6501), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I969 (.Y(N5939), .A0(N6273), .A1(N6487), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I970 (.Y(N6102), .A0(N6273), .A1(N6490), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I971 (.Y(N6253), .A0(N6273), .A1(N6501), .B0(N6411), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I972 (.Y(N6405), .A(N6273), .B(N6411));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I973 (.Y(N5912), .A0(N6273), .A1(N6011), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I974 (.Y(N6081), .A0(N6273), .A1(N6021), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I975 (.Y(N6228), .A0(N6273), .A1(N6501), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I976 (.Y(N6381), .A0(N6273), .A1(N6238), .B0(N6328), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I977 (.Y(N6532), .A0(N6273), .A1(N5877), .B0(N6139), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I978 (.Y(N5978), .A(N6273), .B(N6501));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I979 (.Y(N6275), .A0(N6273), .A1(N6198), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I980 (.Y(N6575), .A0(N6273), .A1(N5877), .B0(inst_cellmath__61[18]), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I981 (.Y(N6183), .A(N6238), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I982 (.Y(N6485), .A0(N6273), .A1(N6411), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I983 (.Y(N6359), .A0(N6273), .A1(N6011), .B0(N6411), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I984 (.Y(N6504), .A(N6273), .B(inst_cellmath__61[18]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I985 (.Y(N6099), .A(N6349), .B(inst_cellmath__61[18]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I986 (.Y(N6544), .A0(N6273), .A1(N6328), .B0(N6487), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I987 (.Y(N5992), .A(N6273), .B(N5877));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I988 (.Y(N6450), .A0(N6273), .A1(N6411), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I989 (.Y(N5894), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I990 (.Y(N6402), .A0(N6273), .A1(N6198), .B0(N6411), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I991 (.Y(N6214), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6328), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I992 (.Y(N6005), .A(N6273), .B(N6238));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I993 (.Y(N6315), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I994 (.Y(N6278), .A0(N6273), .A1(N6241), .B0(N6011), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I995 (.Y(N6186), .A(N6328), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I996 (.Y(N6489), .A0(N6273), .A1(N6198), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I997 (.Y(N5937), .A0(N6273), .A1(N6238), .B0(N6411), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I998 (.Y(N6101), .A(N6273), .B(N6490));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I999 (.Y(N6007), .A0(N6273), .A1(N6490), .B0(N6328), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1000 (.Y(N6461), .A0(N6273), .A1(N6238), .B0(N6241), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1001 (.Y(N6077), .A(N6273), .B(N6198));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1002 (.Y(N6529), .A0(N6273), .A1(N6198), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1003 (.Y(N5974), .A0(N6273), .A1(N6238), .B0(N6501), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1004 (.Y(N6134), .A(N6349), .B(N6011));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1005 (.Y(N5878), .A(N6349), .B(N6241));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1006 (.Y(N5906), .A(N6349), .B(N6501));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1007 (.Y(N6224), .A(N6198), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1008 (.Y(N6459), .A0(N6273), .A1(N5877), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1009 (.Y(N5907), .A0(N6273), .A1(N5877), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1010 (.Y(N6075), .A0(N6273), .A1(N6198), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1011 (.Y(N6225), .A0(N6273), .A1(N5877), .B0(N6411), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1012 (.Y(N6377), .A(N6139), .B(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1013 (.Y(N6527), .A(N6349), .B(N5877));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1014 (.Y(N6132), .A0(N6273), .A1(N6198), .B0(N6238), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1015 (.Y(N6351), .A(N6349), .B(N6328));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1016 (.Y(N6433), .A0(N6273), .A1(N6021), .B0(N6011), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1017 (.Y(N6261), .A(N6241));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1018 (.Y(N6408), .A0(N6273), .A1(N6021), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1019 (.Y(N6560), .A0(N6273), .A1(N6139), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1020 (.Y(N6016), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1021 (.Y(N6168), .A0(N6273), .A1(N6241), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1022 (.Y(N6044), .A0(N6273), .A1(N6198), .B0(N6139), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1023 (.Y(N6350), .A(N6349), .B(N6198));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1024 (.Y(N5945), .A(N6273), .B(N6238));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1025 (.Y(N5887), .A0(N6273), .A1(N6411), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1026 (.Y(N6055), .A0(N6273), .A1(N6487), .B0(N6411), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1027 (.Y(N6260), .A0(N6273), .A1(N6501), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1028 (.Y(N6511), .A0(N6273), .A1(N5877), .B0(N6198), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1029 (.Y(N5954), .A(N6490));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1030 (.Y(N6030), .A0(N6273), .A1(N6487), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1031 (.Y(N6179), .A0(N6273), .A1(N6490), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1032 (.Y(N6337), .A0(N6273), .A1(N6487), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1033 (.Y(N5931), .A0(N6273), .A1(N6411), .B0(N6501), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1034 (.Y(N6167), .A(N6273), .B(N6411));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1035 (.Y(N6070), .A0(N6273), .A1(N6198), .B0(N6021), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1036 (.Y(N6374), .A(N6273), .B(inst_cellmath__61[18]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1037 (.Y(N6129), .A(N6490), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1038 (.Y(N6429), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6241), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1039 (.Y(N6471), .A(inst_cellmath__61[18]), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1040 (.Y(N6193), .A0(N6273), .A1(N6487), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1041 (.Y(N6346), .A0(N6273), .A1(N6238), .B0(N6011), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1042 (.Y(N5942), .A(N6273), .B(N6198));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1043 (.Y(N6255), .A(N6273), .B(N6021));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1044 (.Y(N6012), .A(N6273), .B(N5877));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1045 (.Y(N6466), .A0(N6273), .A1(N6241), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1046 (.Y(N5915), .A0(N6273), .A1(N6501), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1047 (.Y(N6293), .A0(N6273), .A1(N6139), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1048 (.Y(N6440), .A0(N6273), .A1(N5877), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1049 (.Y(N6087), .A0(N6273), .A1(N6490), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1050 (.Y(N6507), .A0(N6273), .A1(N6487), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1051 (.Y(N5952), .A0(N6273), .A1(N6139), .B0(inst_cellmath__61[18]), .B1(N6349));
XNOR2X4 inst_cellmath__195__80__2WWMM_2WWMM_I8329 (.Y(N5911), .A(N704), .B(N5817));
CLKINVX4 inst_cellmath__195__80__2WWMM_2WWMM_I1054 (.Y(N6064), .A(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1055 (.Y(N6244), .A0(N6064), .A1(N6492), .B0(N5928), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1056 (.Y(N6394), .A0(N6064), .A1(inst_cellmath__61[18]), .B0(N6094), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1057 (.Y(N6546), .A0(N6064), .A1(N6224), .B0(N6147), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1058 (.Y(N5994), .A0(N6064), .A1(N6459), .B0(N5996), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1059 (.Y(N6152), .A0(N6064), .A1(N5907), .B0(N6154), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1061 (.Y(N6307), .A0(N6064), .A1(N6075), .B0(N6448), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1062 (.Y(N6452), .A0(N6064), .A1(N6225), .B0(N5898), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1063 (.Y(N5896), .A0(N6064), .A1(N6377), .B0(N6059), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1064 (.Y(N6065), .A0(N6064), .A1(N6527), .B0(N6218), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1065 (.Y(N6216), .A0(N6064), .A1(N6147), .B0(N6370), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1066 (.Y(N6368), .A0(N6064), .A1(N6132), .B0(N5966), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1067 (.Y(N6518), .A0(N6064), .A1(N6351), .B0(N6365), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1068 (.Y(N5964), .A0(N6064), .A1(N6433), .B0(N6281), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1069 (.Y(N6124), .A0(N6064), .A1(N6261), .B0(N5959), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1070 (.Y(N6279), .A0(N6064), .A1(N6408), .B0(N6343), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1071 (.Y(N6426), .A0(N6064), .A1(N6560), .B0(N6492), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1072 (.Y(N6579), .A0(N6064), .A1(N6016), .B0(N5939), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1073 (.Y(N6038), .A0(N6064), .A1(N6168), .B0(N6102), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1074 (.Y(N6188), .A0(N6064), .A1(N6044), .B0(N6253), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1075 (.Y(N6342), .A0(N6064), .A1(N6350), .B0(N6405), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1076 (.Y(N6491), .A(N5911), .B(N5945));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1077 (.Y(N6163), .A0(N6064), .A1(N5906), .B0(N6059), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1078 (.Y(N6318), .A0(N6064), .A1(N5887), .B0(N5912), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1079 (.Y(N6463), .A0(N6064), .A1(N6055), .B0(N6081), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1080 (.Y(N5910), .A0(N6064), .A1(N6275), .B0(N6228), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1081 (.Y(N6079), .A0(N6064), .A1(N6260), .B0(N6381), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1082 (.Y(N6227), .A0(N6064), .A1(N6511), .B0(N6532), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1083 (.Y(N6380), .A0(N6064), .A1(N6315), .B0(N5978), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1084 (.Y(N6531), .A0(N6064), .A1(N5954), .B0(N6275), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1085 (.Y(N5977), .A0(N6064), .A1(N6016), .B0(N6575), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1086 (.Y(N6136), .A0(N6064), .A1(N6349), .B0(N6183), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1087 (.Y(N6290), .A0(N6064), .A1(N6030), .B0(N6485), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1088 (.Y(N6437), .A0(N6064), .A1(N6179), .B0(N6359), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1089 (.Y(N5881), .A0(N6064), .A1(N6337), .B0(N6504), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1090 (.Y(N6048), .A0(N6064), .A1(N5954), .B0(N6099), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1091 (.Y(N6201), .A0(N6064), .A1(N5931), .B0(N5959), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1092 (.Y(N6358), .A(N5911), .B(N6167));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1093 (.Y(N6331), .A0(N6064), .A1(N6070), .B0(N6544), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1094 (.Y(N6476), .A0(N6064), .A1(N6214), .B0(N5992), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1095 (.Y(N5925), .A0(N6064), .A1(N6374), .B0(N6450), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1096 (.Y(N6091), .A0(N6064), .A1(N6129), .B0(N5894), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1097 (.Y(N6242), .A0(N6064), .A1(N6429), .B0(N6402), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1098 (.Y(N6392), .A0(N6064), .A1(N6471), .B0(N6214), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1099 (.Y(N6543), .A0(N6064), .A1(N6193), .B0(N6005), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1100 (.Y(N5991), .A0(N6064), .A1(N6346), .B0(N6315), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1101 (.Y(N6150), .A0(N6064), .A1(N6132), .B0(N6278), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1102 (.Y(N6305), .A0(N6064), .A1(N5942), .B0(N5992), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1103 (.Y(N6449), .A0(N6064), .A1(N6255), .B0(N6186), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1104 (.Y(N5893), .A0(N6064), .A1(N6012), .B0(N6489), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1105 (.Y(N6062), .A0(N6064), .A1(N6260), .B0(N5937), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1106 (.Y(N6213), .A0(N6064), .A1(N6466), .B0(N6101), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1107 (.Y(N6366), .A0(N6064), .A1(N5915), .B0(N6448), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1108 (.Y(N6515), .A0(N6064), .A1(N6351), .B0(N6007), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1109 (.Y(N5961), .A0(N6064), .A1(N6225), .B0(inst_cellmath__61[18]), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1110 (.Y(N6122), .A0(N6064), .A1(N6044), .B0(N6461), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1111 (.Y(N6277), .A0(N6064), .A1(N6381), .B0(N6365), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1112 (.Y(N6424), .A0(N6064), .A1(N6293), .B0(N6077), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1113 (.Y(N6577), .A0(N6064), .A1(N6440), .B0(N6529), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1114 (.Y(N6036), .A0(N6064), .A1(inst_cellmath__61[18]), .B0(N5974), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1115 (.Y(N6185), .A0(N6064), .A1(N6560), .B0(N6134), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1116 (.Y(N6341), .A0(N6064), .A1(N6087), .B0(N5878), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1117 (.Y(N6488), .A0(N6064), .A1(N6507), .B0(N5906), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1118 (.Y(N5936), .A(N6064), .B(N5952));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1119 (.Y(N6251), .A(N6064), .B(N6099));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1120 (.Y(N6146), .A0(N6273), .A1(N6241), .B0(N6411), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1121 (.Y(N6301), .A0(N6273), .A1(N6487), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1122 (.Y(N6447), .A0(N6273), .A1(N6238), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1123 (.Y(N5891), .A0(N6273), .A1(N6198), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1124 (.Y(N6058), .A0(N6273), .A1(N6241), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1125 (.Y(N6210), .A0(N6273), .A1(N6021), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1126 (.Y(N6513), .A0(N6273), .A1(N6198), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1127 (.Y(N5958), .A0(N6273), .A1(N6011), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1128 (.Y(N6120), .A0(N6273), .A1(N6490), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1129 (.Y(N6274), .A0(N6273), .A1(N6501), .B0(N6328), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1130 (.Y(N6422), .A(N6273), .B(N6501));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1131 (.Y(N6182), .A(N6273), .B(inst_cellmath__61[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1132 (.Y(N6389), .A0(N6273), .A1(N6238), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1133 (.Y(N6400), .A0(N6273), .A1(N6011), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1134 (.Y(N6553), .A0(N6273), .A1(N6139), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1135 (.Y(N6526), .A0(N6273), .A1(N6011), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1136 (.Y(N5972), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6011), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1137 (.Y(N6432), .A(N6273), .B(N6490));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1138 (.Y(N6043), .A0(N6273), .A1(N6139), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1139 (.Y(N6259), .A0(N6273), .A1(N6241), .B0(N6021), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1140 (.Y(N6015), .A(N6273), .B(N6241));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1141 (.Y(N6387), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1142 (.Y(N5998), .A0(N6273), .A1(N6021), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1143 (.Y(N6310), .A0(N6273), .A1(N5877), .B0(N6328), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1144 (.Y(N5900), .A0(N6273), .A1(N6487), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1145 (.Y(N6521), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1146 (.Y(N5985), .A0(N6273), .A1(N6328), .B0(N6238), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1147 (.Y(N6127), .A(N6349), .B(N6021));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1148 (.Y(N6581), .A0(N6273), .A1(N6139), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1149 (.Y(N6191), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1150 (.Y(N6344), .A0(N6273), .A1(N6139), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1151 (.Y(N6494), .A0(N6273), .A1(N6490), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1152 (.Y(N5941), .A0(N6273), .A1(N6411), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1153 (.Y(N6104), .A0(N6273), .A1(N6011), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1154 (.Y(N6578), .A0(N6273), .A1(N6411), .B0(inst_cellmath__61[18]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1155 (.Y(N6037), .A0(N6273), .A1(N6198), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1156 (.Y(N5938), .A0(N6273), .A1(N6490), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1157 (.Y(N6404), .A0(N6273), .A1(N6490), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1158 (.Y(N6174), .A0(N6273), .A1(N6021), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1159 (.Y(N6330), .A0(N6273), .A1(N5877), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1160 (.Y(N5923), .A0(N6273), .A1(N6501), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1161 (.Y(N6240), .A0(N6273), .A1(N6328), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1162 (.Y(N6297), .A0(N6273), .A1(N5877), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1163 (.Y(N6541), .A0(N6273), .A1(N6487), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1164 (.Y(N5990), .A0(N6273), .A1(N6011), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1165 (.Y(N6148), .A0(N6273), .A1(N6328), .B0(N6411), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1166 (.Y(N6303), .A0(N6273), .A1(N6139), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1167 (.Y(N6060), .A0(N6273), .A1(N6241), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1168 (.Y(N6211), .A0(N6273), .A1(N6487), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1169 (.Y(N5886), .A0(N6273), .A1(N6238), .B0(N6198), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1170 (.Y(N6460), .A0(N6273), .A1(N6021), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1171 (.Y(N5908), .A0(N6273), .A1(N6238), .B0(N6490), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1172 (.Y(N6206), .A(N5877), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1173 (.Y(N6354), .A0(N6273), .A1(N6490), .B0(N6411), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1174 (.Y(N6264), .A(N6349), .B(N6411));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1175 (.Y(N6510), .A0(N6273), .A1(N6241), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1176 (.Y(N6119), .A0(N6064), .A1(N6055), .B0(N6146), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1177 (.Y(N6272), .A0(N6064), .A1(N6578), .B0(N6301), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1178 (.Y(N6421), .A0(N6064), .A1(N6037), .B0(N6447), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1179 (.Y(N6574), .A0(N6064), .A1(N6087), .B0(N5891), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1180 (.Y(N6033), .A(N6064), .B(N6058));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1181 (.Y(N6483), .A0(N6064), .A1(N6529), .B0(N6210), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1182 (.Y(N5934), .A0(N6064), .A1(N5938), .B0(N6087), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1183 (.Y(N6098), .A(N6513), .B(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1184 (.Y(N6399), .A0(N6064), .A1(N6404), .B0(N5958), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1185 (.Y(N6552), .A0(N6064), .A1(N5958), .B0(N6120), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1186 (.Y(N6002), .A0(N6064), .A1(N6011), .B0(N6274), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1187 (.Y(N6160), .A0(N6064), .A1(N6544), .B0(N6422), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1188 (.Y(N6314), .A0(N6064), .A1(N5900), .B0(N6182), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1189 (.Y(N6458), .A0(N6064), .A1(N6527), .B0(N6278), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1190 (.Y(N5904), .A0(N6064), .A1(N6099), .B0(N6389), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1191 (.Y(N6074), .A(N6064), .B(N6471));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1192 (.Y(N6525), .A0(N6064), .A1(inst_cellmath__61[17]), .B0(N6400), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1193 (.Y(N5971), .A0(N6064), .A1(inst_cellmath__61[18]), .B0(N6553), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1194 (.Y(N6131), .A0(N6064), .A1(N6273), .B0(N6183), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1195 (.Y(N6285), .A0(N6064), .A1(N6273), .B0(N6349), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1196 (.Y(N6431), .A(N6064), .B(N6273));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1197 (.Y(N6042), .A(N5911), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1198 (.Y(N6107), .A0(N6064), .A1(N6174), .B0(N6526), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1199 (.Y(N6258), .A0(N6064), .A1(N6330), .B0(N5972), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1200 (.Y(N6559), .A(N5911), .B(N5923));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1201 (.Y(N6325), .A0(N6064), .A1(N5915), .B0(N6432), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1202 (.Y(N6469), .A0(N6064), .A1(N6240), .B0(N6043), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1203 (.Y(N5918), .A0(N6064), .A1(N6297), .B0(N6527), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1204 (.Y(N6086), .A0(N6064), .A1(N6541), .B0(N6365), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1205 (.Y(N6234), .A0(N6064), .A1(N5990), .B0(N6408), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1206 (.Y(N6386), .A0(N6064), .A1(N6148), .B0(N6259), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1207 (.Y(N6537), .A0(N6064), .A1(N6303), .B0(N6186), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1208 (.Y(N5983), .A0(N6064), .A1(N6400), .B0(N6015), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1209 (.Y(N6140), .A0(N6064), .A1(N6387), .B0(N6167), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1210 (.Y(N6295), .A0(N6064), .A1(N6060), .B0(N6526), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1211 (.Y(N6442), .A0(N6064), .A1(N6211), .B0(N6387), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1212 (.Y(N5884), .A0(N6064), .A1(N5886), .B0(N6293), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1213 (.Y(N6053), .A0(N6064), .A1(N6224), .B0(N6005), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1214 (.Y(N6115), .A(N5911), .B(N6005));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1215 (.Y(N6570), .A0(N6064), .A1(N6504), .B0(N6402), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1216 (.Y(N6027), .A0(N6064), .A1(N6422), .B0(N6432), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1217 (.Y(N6177), .A0(N6064), .A1(N6492), .B0(N6349), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1218 (.Y(N6334), .A(N6064), .B(N6030));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1219 (.Y(N5929), .A0(N6064), .A1(N6365), .B0(N5959), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1220 (.Y(N6095), .A0(N6064), .A1(N6303), .B0(N6281), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1221 (.Y(N6246), .A0(N6064), .A1(N6460), .B0(N5906), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1222 (.Y(N6396), .A0(N6064), .A1(N5908), .B0(N5998), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1223 (.Y(N6548), .A0(N6064), .A1(N6460), .B0(N6485), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1224 (.Y(N5997), .A0(N6064), .A1(N6575), .B0(N6310), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1225 (.Y(N6155), .A0(N6064), .A1(N6330), .B0(N6433), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1226 (.Y(N6309), .A0(N6064), .A1(N6447), .B0(N5900), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1227 (.Y(N6454), .A0(N6064), .A1(N6408), .B0(N5937), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1228 (.Y(N5899), .A0(N6064), .A1(N6206), .B0(N6485), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1229 (.Y(N6068), .A0(N6064), .A1(N6102), .B0(N6218), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1230 (.Y(N6219), .A0(N6064), .A1(N6005), .B0(N6521), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1231 (.Y(N6371), .A0(N6064), .A1(N6354), .B0(N5985), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1232 (.Y(N6520), .A0(N6064), .A1(N6281), .B0(N6127), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1233 (.Y(N5967), .A0(N6064), .A1(N6264), .B0(N6581), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1234 (.Y(N6126), .A0(N6064), .A1(N6510), .B0(N6343), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1235 (.Y(N6282), .A0(N6064), .A1(N5972), .B0(N6191), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1236 (.Y(N6427), .A0(N6064), .A1(N6260), .B0(N6344), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1237 (.Y(N6580), .A(N6494), .B(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1238 (.Y(N6189), .A(N5941), .B(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1239 (.Y(N6493), .A0(N6064), .A1(inst_cellmath__61[17]), .B0(N6104), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1240 (.Y(N5940), .A0(N6064), .A1(N5954), .B0(N6448), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1241 (.Y(N6103), .A0(N6064), .A1(N5886), .B0(N5945), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1242 (.Y(N6254), .A0(N6064), .A1(N5945), .B0(N6350), .B1(N5911));
XNOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8330 (.Y(N5962), .A(N5817), .B(N705));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1245 (.Y(N5989), .A(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1246 (.Y(N6320), .A0(N5989), .A1(N6119), .B0(N6244), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1247 (.Y(N6464), .A0(N5989), .A1(N6272), .B0(N6394), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1248 (.Y(N5913), .A0(N5989), .A1(N6421), .B0(N6546), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1249 (.Y(N6082), .A0(N5989), .A1(N6574), .B0(N5994), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1250 (.Y(N6229), .A0(N5989), .A1(N6033), .B0(N6152), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1251 (.Y(N6382), .A0(N5989), .A1(N6483), .B0(N6307), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1252 (.Y(N6533), .A0(N5989), .A1(N5934), .B0(N6452), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1253 (.Y(N5979), .A0(N5989), .A1(N6098), .B0(N5896), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1254 (.Y(N6137), .A0(N5989), .A1(N6399), .B0(N6065), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1255 (.Y(N6291), .A0(N5989), .A1(N6552), .B0(N6216), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1256 (.Y(N6438), .A0(N5989), .A1(N6002), .B0(N6368), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1257 (.Y(N5882), .A0(N5989), .A1(N6160), .B0(N6518), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1258 (.Y(N6049), .A0(N5989), .A1(N6314), .B0(N5964), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1259 (.Y(N6202), .A0(N5989), .A1(N6458), .B0(N6124), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1260 (.Y(N6360), .A0(N5989), .A1(N5904), .B0(N6279), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1261 (.Y(N6505), .A0(N5989), .A1(N6074), .B0(N6426), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1262 (.Y(N5950), .A0(N5989), .A1(N6525), .B0(N6579), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1263 (.Y(N6112), .A0(N5989), .A1(N5971), .B0(N6038), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1264 (.Y(N6267), .A0(N5989), .A1(N6131), .B0(N6188), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1265 (.Y(N6414), .A0(N5989), .A1(N6285), .B0(N6342), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1266 (.Y(N6566), .A0(N5989), .A1(N6431), .B0(N6491), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1267 (.Y(N6477), .A0(N5989), .A1(N6107), .B0(N6163), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1268 (.Y(N5926), .A0(N5989), .A1(N6258), .B0(N6318), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1269 (.Y(N6092), .A0(N5989), .A1(N6227), .B0(N6463), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1270 (.Y(N6243), .A0(N5989), .A1(N6559), .B0(N5910), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1271 (.Y(N6393), .A0(N5989), .A1(N6325), .B0(N6079), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1272 (.Y(N6545), .A0(N5989), .A1(N6469), .B0(N6227), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1273 (.Y(N5993), .A0(N5989), .A1(N5918), .B0(N6380), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1274 (.Y(N6151), .A0(N5989), .A1(N6086), .B0(N6531), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1275 (.Y(N6306), .A0(N5989), .A1(N6234), .B0(N5977), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1276 (.Y(N6451), .A0(N5989), .A1(N6386), .B0(N6136), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1277 (.Y(N5895), .A0(N5989), .A1(N6537), .B0(N6290), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1278 (.Y(N6063), .A0(N5989), .A1(N5983), .B0(N6437), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1279 (.Y(N6215), .A0(N5989), .A1(N6140), .B0(N5881), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1280 (.Y(N6367), .A0(N5989), .A1(N6295), .B0(N6048), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1281 (.Y(N6516), .A0(N5989), .A1(N6442), .B0(N6201), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1282 (.Y(N5963), .A0(N5989), .A1(N5884), .B0(N6358), .B1(N5962));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1283 (.Y(N6123), .A(N5989), .B(N6053));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1284 (.Y(N5975), .A(N6064), .B(N6224));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1285 (.Y(N6425), .A(N5962), .B(N5975));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1286 (.Y(N6252), .A0(N5989), .A1(N6570), .B0(N6331), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1287 (.Y(N6403), .A0(N5989), .A1(N6027), .B0(N6476), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1288 (.Y(N6555), .A0(N5989), .A1(N6177), .B0(N5925), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1289 (.Y(N6008), .A0(N5989), .A1(N6334), .B0(N6091), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1290 (.Y(N6162), .A0(N5989), .A1(N5929), .B0(N6242), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1291 (.Y(N6317), .A0(N5989), .A1(N6095), .B0(N6392), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1292 (.Y(N6462), .A0(N5989), .A1(N6246), .B0(N6543), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1293 (.Y(N5909), .A0(N5989), .A1(N6396), .B0(N5991), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1294 (.Y(N6078), .A0(N5989), .A1(N6548), .B0(N6150), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1295 (.Y(N6226), .A0(N5989), .A1(N5997), .B0(N6305), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1296 (.Y(N6379), .A0(N5989), .A1(N6155), .B0(N6449), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1297 (.Y(N6530), .A0(N5989), .A1(N6309), .B0(N5893), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1298 (.Y(N5976), .A0(N5989), .A1(N6454), .B0(N6062), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1299 (.Y(N6135), .A0(N5989), .A1(N5899), .B0(N6213), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1300 (.Y(N6288), .A0(N5989), .A1(N6068), .B0(N6366), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1301 (.Y(N6435), .A0(N5989), .A1(N6219), .B0(N6515), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1302 (.Y(N5879), .A0(N5989), .A1(N6371), .B0(N5961), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1303 (.Y(N6046), .A0(N5989), .A1(N6520), .B0(N6122), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1304 (.Y(N6199), .A0(N5989), .A1(N5967), .B0(N6277), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1305 (.Y(N6356), .A0(N5989), .A1(N6126), .B0(N6424), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1306 (.Y(N6502), .A0(N5989), .A1(N6282), .B0(N6577), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1307 (.Y(N5948), .A0(N5989), .A1(N6427), .B0(N6036), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1308 (.Y(N6110), .A0(N5989), .A1(N6580), .B0(N6185), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1309 (.Y(N6265), .A0(N5989), .A1(N6189), .B0(N6341), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1310 (.Y(N6412), .A0(N5989), .A1(N6493), .B0(N6488), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1311 (.Y(N6564), .A0(N5989), .A1(N5940), .B0(N5936), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1312 (.Y(N6022), .A0(N5989), .A1(N6103), .B0(N6251), .B1(N5962));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1313 (.Y(N6172), .A(N5962), .B(N6254));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1314 (.Y(N6355), .A(N6064), .B(N6350));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1315 (.Y(N5921), .A(N5962), .B(N6355));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1316 (.Y(N6561), .A0(N6273), .A1(N6501), .B0(N5877), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1317 (.Y(N6472), .A(N6349), .B(N6238));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1318 (.Y(N5986), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1319 (.Y(N6298), .A0(N6273), .A1(N6487), .B0(N6328), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1320 (.Y(N6444), .A(N6487));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1321 (.Y(N5888), .A0(N6273), .A1(N6411), .B0(N6328), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1322 (.Y(N6056), .A0(N6273), .A1(N5877), .B0(N6501), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1323 (.Y(N6207), .A0(N6273), .A1(N6241), .B0(inst_cellmath__61[17]), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1324 (.Y(N6071), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1325 (.Y(N6221), .A0(N6273), .A1(N6238), .B0(inst_cellmath__61[17]), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1326 (.Y(N6322), .A(N6349), .B(inst_cellmath__61[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1327 (.Y(N6231), .A0(N6273), .A1(N6411), .B0(N6011), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1328 (.Y(N6294), .A0(N6273), .A1(N6011), .B0(N6238), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1329 (.Y(N6441), .A0(N6273), .A1(N6487), .B0(inst_cellmath__61[18]), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1330 (.Y(N6051), .A(N6411), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1331 (.Y(N6568), .A0(N6273), .A1(N6411), .B0(N6021), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1332 (.Y(N6025), .A(N6273), .B(N6011));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1333 (.Y(N6479), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N5877), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1334 (.Y(N6117), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6021), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1335 (.Y(N6066), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6490), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1336 (.Y(N6076), .A(N6273), .B(N6487));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1337 (.Y(N6019), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6411), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1338 (.Y(N6237), .A(N6238));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1339 (.Y(N6391), .A0(N6273), .A1(N6490), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1340 (.Y(N5988), .A0(N6273), .A1(N6241), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1341 (.Y(N6302), .A0(N6273), .A1(N6241), .B0(N6328), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1342 (.Y(N6034), .A0(N6273), .A1(N5877), .B0(N6238), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1343 (.Y(N6484), .A(N6501));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1344 (.Y(N6401), .A0(N6273), .A1(N6328), .B0(N6241), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1345 (.Y(N6004), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6139), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1346 (.Y(N5905), .A0(N6273), .A1(N6238), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1347 (.Y(N6286), .A0(N6273), .A1(N6139), .B0(N6241), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1348 (.Y(N6470), .A(N6501), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1349 (.Y(N6235), .A0(N6064), .A1(N5941), .B0(N6365), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1350 (.Y(N6388), .A0(N6064), .A1(N6261), .B0(N5878), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1351 (.Y(N6538), .A0(N6064), .A1(N6147), .B0(N6005), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1352 (.Y(N5984), .A0(N6064), .A1(N5966), .B0(N6561), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1353 (.Y(N6142), .A0(N6064), .A1(N6206), .B0(N6381), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1354 (.Y(N6296), .A0(N6064), .A1(N6349), .B0(N6532), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1355 (.Y(N6443), .A0(N6064), .A1(N5992), .B0(N6275), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1356 (.Y(N5885), .A0(N6064), .A1(N6349), .B0(N6472), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1357 (.Y(N6054), .A0(N6064), .A1(N6315), .B0(N6273), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1358 (.Y(N6205), .A0(N6064), .A1(N6389), .B0(N6510), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1359 (.Y(N6363), .A0(N6064), .A1(N6489), .B0(N5986), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1360 (.Y(N6509), .A0(N6064), .A1(N6315), .B0(N6191), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1361 (.Y(N5955), .A0(N6064), .A1(N6076), .B0(N6298), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1362 (.Y(N6116), .A0(N6064), .A1(N6221), .B0(N6444), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1363 (.Y(N6270), .A0(N6064), .A1(N6129), .B0(N5888), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1364 (.Y(N6417), .A0(N6064), .A1(N6117), .B0(N6056), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1365 (.Y(N6571), .A0(N6064), .A1(N6102), .B0(N6207), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1366 (.Y(N6028), .A0(N6064), .A1(N5931), .B0(N6275), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1367 (.Y(N6178), .A0(N6064), .A1(N6167), .B0(N6132), .B1(N5911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1368 (.Y(N6335), .A(N5945), .B(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1369 (.Y(N5999), .A0(N6064), .A1(N5931), .B0(N5894), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1370 (.Y(N6156), .A0(N6064), .A1(N6019), .B0(N6344), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1371 (.Y(N6311), .A0(N6064), .A1(N6275), .B0(N6104), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1372 (.Y(N6455), .A0(N6064), .A1(N5886), .B0(N6015), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1373 (.Y(N5901), .A0(N6064), .A1(N6297), .B0(N5996), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1374 (.Y(N6069), .A0(N6064), .A1(N6275), .B0(N6365), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1375 (.Y(N6220), .A0(N6064), .A1(N6561), .B0(N6527), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1376 (.Y(N6373), .A0(N6064), .A1(N6237), .B0(N5959), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1377 (.Y(N6522), .A0(N6064), .A1(N6391), .B0(N6071), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1378 (.Y(N5968), .A0(N6064), .A1(N6404), .B0(N6221), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1379 (.Y(N6128), .A0(N6064), .A1(N5988), .B0(N6260), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1380 (.Y(N6283), .A0(N6064), .A1(N6400), .B0(N6578), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1381 (.Y(N6428), .A0(N6064), .A1(N6302), .B0(N6011), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1382 (.Y(N6582), .A0(N6064), .A1(N6253), .B0(inst_cellmath__61[18]), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1383 (.Y(N6039), .A0(N6064), .A1(N6117), .B0(N6510), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1384 (.Y(N6192), .A0(N6064), .A1(N6448), .B0(N6402), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1385 (.Y(N6345), .A0(N6064), .A1(N6260), .B0(N6350), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1386 (.Y(N6495), .A0(N6064), .A1(N5906), .B0(N5945), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1387 (.Y(N6556), .A0(N6064), .A1(N6034), .B0(N6132), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1388 (.Y(N6010), .A0(N6064), .A1(N6034), .B0(N6148), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1389 (.Y(N6164), .A0(N6064), .A1(N6060), .B0(N6322), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1390 (.Y(N6321), .A0(N6064), .A1(N6484), .B0(N6575), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1391 (.Y(N6465), .A0(N6064), .A1(N5972), .B0(N6231), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1392 (.Y(N5914), .A0(N6064), .A1(N5959), .B0(N5985), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1393 (.Y(N6083), .A0(N6064), .A1(N6401), .B0(N6448), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1394 (.Y(N6230), .A0(N6064), .A1(N6059), .B0(N5942), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1395 (.Y(N6383), .A0(N6064), .A1(N6004), .B0(N6294), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1396 (.Y(N6534), .A0(N6064), .A1(N5898), .B0(N6441), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1397 (.Y(N5980), .A0(N6064), .A1(N5942), .B0(N6330), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1398 (.Y(N6138), .A0(N6064), .A1(N5905), .B0(N6051), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1399 (.Y(N6292), .A0(N6064), .A1(N6037), .B0(N6374), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1400 (.Y(N6439), .A0(N6064), .A1(N6510), .B0(N6374), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1401 (.Y(N5883), .A0(N6064), .A1(N5923), .B0(N6568), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1402 (.Y(N6050), .A0(N6064), .A1(N6056), .B0(N6025), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1403 (.Y(N6203), .A0(N6064), .A1(N6060), .B0(N6479), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1404 (.Y(N6361), .A0(N6064), .A1(N6389), .B0(N6471), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1405 (.Y(N6506), .A0(N6064), .A1(N6286), .B0(N6030), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1406 (.Y(N5951), .A0(N6064), .A1(N6044), .B0(N6117), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1407 (.Y(N6113), .A0(N6064), .A1(N5985), .B0(N6211), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1408 (.Y(N6268), .A0(N6064), .A1(N6337), .B0(N6444), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1409 (.Y(N6415), .A0(N6064), .A1(N6275), .B0(N6561), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1410 (.Y(N6567), .A0(N6064), .A1(N6310), .B0(N6139), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1411 (.Y(N6024), .A0(N6064), .A1(N6259), .B0(N6016), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1412 (.Y(N6175), .A0(N6064), .A1(N6440), .B0(N6066), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1413 (.Y(N6332), .A0(N6064), .A1(N6019), .B0(N6077), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1414 (.Y(N6478), .A0(N6064), .A1(N6167), .B0(N6273), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1415 (.Y(N6418), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6021), .B1(N6349));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1416 (.Y(N5924), .A(N6273), .B(N6487));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1417 (.Y(N6542), .A0(N6273), .A1(N6501), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1418 (.Y(N6149), .A0(N6273), .A1(N6011), .B0(N6328), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1419 (.Y(N6304), .A(N6021));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1420 (.Y(N5892), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6411), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1421 (.Y(N6061), .A0(N6273), .A1(N6490), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1422 (.Y(N6212), .A0(N6273), .A1(N6411), .B0(N6238), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1423 (.Y(N6145), .A(N5877));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1424 (.Y(N5957), .A(N6273), .B(inst_cellmath__61[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1425 (.Y(N6003), .A0(N6273), .A1(N6139), .B0(N6501), .B1(N6349));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1426 (.Y(N6141), .A(N6198));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1427 (.Y(N6372), .A(N6021), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1428 (.Y(N6190), .A0(N6273), .A1(N6198), .B0(N6490), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1429 (.Y(N6009), .A0(N6273), .A1(inst_cellmath__61[17]), .B0(N6490), .B1(N6349));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1430 (.Y(N6517), .A(N6487), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1431 (.Y(N6187), .A0(N6273), .A1(inst_cellmath__61[18]), .B0(N6487), .B1(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1432 (.Y(N6289), .A0(N6064), .A1(N5990), .B0(N6255), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1433 (.Y(N6436), .A0(N6064), .A1(N6070), .B0(N6578), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1434 (.Y(N5880), .A0(N6064), .A1(N6141), .B0(N6076), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1435 (.Y(N6047), .A0(N6064), .A1(N6206), .B0(N6418), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1436 (.Y(N6200), .A0(N6064), .A1(N6186), .B0(N6485), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1437 (.Y(N6357), .A0(N6064), .A1(N6206), .B0(N6231), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1438 (.Y(N6503), .A0(N6064), .A1(N6302), .B0(N6127), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1439 (.Y(N5949), .A0(N6064), .A1(N6104), .B0(N5924), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1440 (.Y(N6111), .A0(N6064), .A1(N6354), .B0(N6056), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1441 (.Y(N6266), .A0(N6064), .A1(N6221), .B0(N6542), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1442 (.Y(N6413), .A0(N6064), .A1(N6044), .B0(N5939), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1443 (.Y(N6565), .A0(N6064), .A1(N6087), .B0(N6149), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1444 (.Y(N6023), .A0(N6064), .A1(N5892), .B0(N6304), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1445 (.Y(N6173), .A0(N6064), .A1(N6007), .B0(N6286), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1446 (.Y(N6329), .A0(N6064), .A1(N5941), .B0(N5892), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1447 (.Y(N6475), .A0(N6064), .A1(N6183), .B0(N6061), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1448 (.Y(N5922), .A0(N6064), .A1(N6273), .B0(N6212), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1449 (.Y(N6090), .A0(N6064), .A1(N6349), .B0(N6273), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1450 (.Y(N6239), .A(N6064), .B(N6273));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1451 (.Y(N6514), .A0(N6064), .A1(N6372), .B0(N6297), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1452 (.Y(N5960), .A0(N6064), .A1(N5978), .B0(N5985), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1453 (.Y(N6121), .A0(N6064), .A1(N6051), .B0(N6389), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1454 (.Y(N6276), .A0(N6064), .A1(N5891), .B0(N6418), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1455 (.Y(N6423), .A0(N6064), .A1(N5928), .B0(N6553), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1456 (.Y(N6576), .A0(N6064), .A1(N6190), .B0(N6581), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1457 (.Y(N6035), .A0(N6064), .A1(N6206), .B0(N6275), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1458 (.Y(N6184), .A0(N6064), .A1(N6273), .B0(N5888), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1459 (.Y(N6340), .A0(N6064), .A1(N5924), .B0(N6471), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1460 (.Y(N6486), .A0(N6064), .A1(N6009), .B0(N6129), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1461 (.Y(N5935), .A0(N6064), .A1(N6418), .B0(N6149), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1462 (.Y(N6100), .A0(N6064), .A1(N6183), .B0(N5954), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1463 (.Y(N6250), .A0(N6064), .A1(N6224), .B0(N5886), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1464 (.Y(N6006), .A0(N6064), .A1(inst_cellmath__61[17]), .B0(N5996), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1465 (.Y(N6161), .A0(N6064), .A1(inst_cellmath__61[18]), .B0(N6043), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1466 (.Y(N6316), .A0(N6064), .A1(N6349), .B0(N6167), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1467 (.Y(N6378), .A0(N6064), .A1(N6484), .B0(N6298), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1468 (.Y(N6528), .A0(N6064), .A1(N6542), .B0(N6147), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1469 (.Y(N5973), .A0(N6064), .A1(N6087), .B0(N6418), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1470 (.Y(N6133), .A0(N6064), .A1(N6448), .B0(N6418), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1471 (.Y(N6287), .A0(N6064), .A1(N6231), .B0(N6441), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1472 (.Y(N6434), .A0(N6064), .A1(N6459), .B0(N6191), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1473 (.Y(N5876), .A0(N6064), .A1(N6127), .B0(N6034), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1474 (.Y(N6045), .A0(N6064), .A1(N5886), .B0(N6297), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1475 (.Y(N6197), .A0(N6064), .A1(N6433), .B0(N6575), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1476 (.Y(N6352), .A0(N6064), .A1(N6568), .B0(N6145), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1477 (.Y(N6499), .A0(N6064), .A1(N6077), .B0(N6117), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1478 (.Y(N5947), .A0(N6064), .A1(N5974), .B0(N6059), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1479 (.Y(N6108), .A0(N6064), .A1(N6190), .B0(inst_cellmath__61[17]), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1480 (.Y(N6262), .A0(N6064), .A1(N6099), .B0(N6404), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1481 (.Y(N6410), .A0(N6064), .A1(N6517), .B0(N6510), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1482 (.Y(N6562), .A0(N6064), .A1(N6099), .B0(N6087), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1483 (.Y(N6017), .A0(N6064), .A1(N6055), .B0(N5957), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1484 (.Y(N6171), .A0(N6064), .A1(N6575), .B0(N6387), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1485 (.Y(N6326), .A0(N6064), .A1(N6187), .B0(N6433), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1486 (.Y(N6474), .A0(N6064), .A1(N6005), .B0(N5938), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1487 (.Y(N5920), .A0(N6064), .A1(N6011), .B0(N6044), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1488 (.Y(N6088), .A(N5911), .B(N6139));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1489 (.Y(N6539), .A(N6064), .B(N6349));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1490 (.Y(N6144), .A0(N6064), .A1(N5958), .B0(N6011), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1491 (.Y(N6299), .A0(N6064), .A1(N6429), .B0(N6261), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1492 (.Y(N6446), .A0(N6064), .A1(N6007), .B0(N6310), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1493 (.Y(N5890), .A0(N6064), .A1(N6402), .B0(N6003), .B1(N5911));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1494 (.Y(N6057), .A0(N6064), .A1(N6470), .B0(N5959), .B1(N5911));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1495 (.Y(N6209), .A(N6064), .B(N6099));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1496 (.Y(N6420), .A0(N5989), .A1(N6289), .B0(N6235), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1497 (.Y(N6573), .A0(N5989), .A1(N6436), .B0(N6388), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1498 (.Y(N6031), .A0(N5989), .A1(N5880), .B0(N6538), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1499 (.Y(N6181), .A0(N5989), .A1(N6047), .B0(N5984), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1500 (.Y(N6339), .A0(N5989), .A1(N6200), .B0(N6142), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1501 (.Y(N6481), .A0(N5989), .A1(N6357), .B0(N6296), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1502 (.Y(N5933), .A0(N5989), .A1(N6503), .B0(N6443), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1503 (.Y(N6096), .A0(N5989), .A1(N5949), .B0(N5885), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1504 (.Y(N6248), .A0(N5989), .A1(N6111), .B0(N6054), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1505 (.Y(N6398), .A0(N5989), .A1(N6266), .B0(N6205), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1506 (.Y(N6550), .A0(N5989), .A1(N6413), .B0(N6363), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1507 (.Y(N6000), .A0(N5989), .A1(N6565), .B0(N6509), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1508 (.Y(N6159), .A0(N5989), .A1(N6023), .B0(N5955), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1509 (.Y(N6312), .A0(N5989), .A1(N6173), .B0(N6116), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1510 (.Y(N6456), .A0(N5989), .A1(N6329), .B0(N6270), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1511 (.Y(N5903), .A0(N5989), .A1(N6475), .B0(N6417), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1512 (.Y(N6072), .A0(N5989), .A1(N5922), .B0(N6571), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1513 (.Y(N6223), .A0(N5989), .A1(N6090), .B0(N6028), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1514 (.Y(N6376), .A0(N5989), .A1(N6239), .B0(N6178), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1515 (.Y(N6523), .A0(N5989), .A1(N6239), .B0(N6335), .B1(N5962));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I1516 (.Y(N5970), .A0N(N6349), .A1N(N5911), .B0(N5989));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1517 (.Y(N6040), .A0(N5989), .A1(N6514), .B0(N5999), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1518 (.Y(N6195), .A0(N5989), .A1(N5960), .B0(N6156), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1519 (.Y(N6348), .A0(N5989), .A1(N6121), .B0(N6311), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1520 (.Y(N6496), .A0(N5989), .A1(N6276), .B0(N6455), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1521 (.Y(N5944), .A0(N5989), .A1(N6423), .B0(N5901), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1522 (.Y(N6106), .A0(N5989), .A1(N6576), .B0(N6069), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1523 (.Y(N6256), .A0(N5989), .A1(N6035), .B0(N6220), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1524 (.Y(N6407), .A0(N5989), .A1(N6184), .B0(N6373), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1525 (.Y(N6558), .A0(N5989), .A1(N6340), .B0(N6522), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1526 (.Y(N6013), .A0(N5989), .A1(N6486), .B0(N5968), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1527 (.Y(N6166), .A0(N5989), .A1(N5935), .B0(N6128), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1528 (.Y(N6324), .A0(N5989), .A1(N6100), .B0(N6283), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1529 (.Y(N6467), .A0(N5989), .A1(N6250), .B0(N6428), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1530 (.Y(N5917), .A0(N5989), .A1(N6335), .B0(N6582), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1531 (.Y(N6085), .A0(N5989), .A1(N6006), .B0(N6039), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1532 (.Y(N6232), .A0(N5989), .A1(N6161), .B0(N6192), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1533 (.Y(N6385), .A0(N5989), .A1(N6316), .B0(N6345), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1534 (.Y(N6536), .A0(N5989), .A1(N6064), .B0(N6495), .B1(N5962));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1535 (.Y(N6020), .A(N5911), .B(N6405));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1536 (.Y(N5981), .A(N6020), .B(N5989));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1537 (.Y(N6052), .A0(N5989), .A1(N6378), .B0(N6556), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1538 (.Y(N6204), .A0(N5989), .A1(N6528), .B0(N6010), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1539 (.Y(N6362), .A0(N5989), .A1(N5973), .B0(N6164), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1540 (.Y(N6508), .A0(N5989), .A1(N6133), .B0(N6321), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1541 (.Y(N5953), .A0(N5989), .A1(N6287), .B0(N6465), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1542 (.Y(N6114), .A0(N5989), .A1(N6434), .B0(N5914), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1543 (.Y(N6269), .A0(N5989), .A1(N5876), .B0(N6083), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1544 (.Y(N6416), .A0(N5989), .A1(N6045), .B0(N6230), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1545 (.Y(N6569), .A0(N5989), .A1(N6197), .B0(N6383), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1546 (.Y(N6026), .A0(N5989), .A1(N6352), .B0(N6534), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1547 (.Y(N6176), .A0(N5989), .A1(N6499), .B0(N5980), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1548 (.Y(N6333), .A0(N5989), .A1(N5947), .B0(N6138), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1549 (.Y(N6480), .A0(N5989), .A1(N6108), .B0(N6292), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1550 (.Y(N5927), .A0(N5989), .A1(N6262), .B0(N6439), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1551 (.Y(N6093), .A0(N5989), .A1(N6410), .B0(N5883), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1552 (.Y(N6245), .A0(N5989), .A1(N6562), .B0(N6050), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1553 (.Y(N6395), .A0(N5989), .A1(N6017), .B0(N6203), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1554 (.Y(N6547), .A0(N5989), .A1(N6171), .B0(N6361), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1555 (.Y(N5995), .A0(N5989), .A1(N6326), .B0(N6506), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1556 (.Y(N6153), .A0(N5989), .A1(N6474), .B0(N5951), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1557 (.Y(N6308), .A0(N5989), .A1(N5920), .B0(N6113), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1558 (.Y(N6453), .A0(N5989), .A1(N6088), .B0(N6268), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1559 (.Y(N5897), .A0(N5989), .A1(N6539), .B0(N6415), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1560 (.Y(N6067), .A0(N5989), .A1(N6144), .B0(N6567), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1561 (.Y(N6217), .A0(N5989), .A1(N6299), .B0(N6024), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1562 (.Y(N6369), .A0(N5989), .A1(N6446), .B0(N6175), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1563 (.Y(N6519), .A0(N5989), .A1(N5890), .B0(N6332), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1564 (.Y(N5965), .A0(N5989), .A1(N6057), .B0(N6478), .B1(N5962));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1565 (.Y(N6125), .A0(N5989), .A1(N6209), .B0(N6358), .B1(N5962));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I1566 (.Y(N6280), .A0N(N6064), .A1N(N6470), .B0(N5962));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1567 (.Y(N6554), .A(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1568 (.Y(N742), .A0(N6554), .A1(N6420), .B0(N6320), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1569 (.Y(N743), .A0(N6554), .A1(N6573), .B0(N6464), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1570 (.Y(N744), .A0(N6554), .A1(N6031), .B0(N5913), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1571 (.Y(N745), .A0(N6554), .A1(N6181), .B0(N6082), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1572 (.Y(N746), .A0(N6554), .A1(N6339), .B0(N6229), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1573 (.Y(N747), .A0(N6554), .A1(N6481), .B0(N6382), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1574 (.Y(N748), .A0(N6554), .A1(N5933), .B0(N6533), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1575 (.Y(N749), .A0(N6554), .A1(N6096), .B0(N5979), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1576 (.Y(N750), .A0(N6554), .A1(N6248), .B0(N6137), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1577 (.Y(N751), .A0(N6554), .A1(N6398), .B0(N6291), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1578 (.Y(N752), .A0(N6554), .A1(N6550), .B0(N6438), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1579 (.Y(N753), .A0(N6554), .A1(N6000), .B0(N5882), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1580 (.Y(N754), .A0(N6554), .A1(N6159), .B0(N6049), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1581 (.Y(N755), .A0(N6554), .A1(N6312), .B0(N6202), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1582 (.Y(N756), .A0(N6554), .A1(N6456), .B0(N6360), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1583 (.Y(N757), .A0(N6554), .A1(N5903), .B0(N6505), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1584 (.Y(N758), .A0(N6554), .A1(N6072), .B0(N5950), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1585 (.Y(N759), .A0(N6554), .A1(N6223), .B0(N6112), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1586 (.Y(N760), .A0(N6554), .A1(N6376), .B0(N6267), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1587 (.Y(N761), .A0(N6554), .A1(N6523), .B0(N6414), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1588 (.Y(N762), .A0(N6554), .A1(N5970), .B0(N6566), .B1(inst_cellmath__61[22]));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I1589 (.Y(N763), .A0N(N5989), .A1N(N6042), .B0(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1590 (.Y(inst_cellmath__197[0]), .A0(N6554), .A1(N6040), .B0(N6477), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1591 (.Y(inst_cellmath__197[1]), .A0(N6554), .A1(N6195), .B0(N5926), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1592 (.Y(inst_cellmath__197[2]), .A0(N6554), .A1(N6348), .B0(N6092), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1593 (.Y(inst_cellmath__197[3]), .A0(N6554), .A1(N6496), .B0(N6243), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1594 (.Y(inst_cellmath__197[4]), .A0(N6554), .A1(N5944), .B0(N6393), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1595 (.Y(inst_cellmath__197[5]), .A0(N6554), .A1(N6106), .B0(N6545), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1596 (.Y(inst_cellmath__197[6]), .A0(N6554), .A1(N6256), .B0(N5993), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1597 (.Y(inst_cellmath__197[7]), .A0(N6554), .A1(N6407), .B0(N6151), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1598 (.Y(inst_cellmath__197[8]), .A0(N6554), .A1(N6558), .B0(N6306), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1599 (.Y(inst_cellmath__197[9]), .A0(N6554), .A1(N6013), .B0(N6451), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1600 (.Y(inst_cellmath__197[10]), .A0(N6554), .A1(N6166), .B0(N5895), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1601 (.Y(inst_cellmath__197[11]), .A0(N6554), .A1(N6324), .B0(N6063), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1602 (.Y(inst_cellmath__197[12]), .A0(N6554), .A1(N6467), .B0(N6215), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1603 (.Y(inst_cellmath__197[13]), .A0(N6554), .A1(N5917), .B0(N6367), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1604 (.Y(inst_cellmath__197[14]), .A0(N6554), .A1(N6085), .B0(N6516), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1605 (.Y(inst_cellmath__197[15]), .A0(N6554), .A1(N6232), .B0(N5963), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1606 (.Y(inst_cellmath__197[16]), .A0(N6554), .A1(N6385), .B0(N6123), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1607 (.Y(inst_cellmath__197[17]), .A0(N6554), .A1(N6536), .B0(N6425), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1608 (.Y(inst_cellmath__197[18]), .A0(N6554), .A1(N5981), .B0(N6425), .B1(inst_cellmath__61[22]));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I1609 (.Y(inst_cellmath__197[19]), .A0N(N5989), .A1N(N6115), .B0(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1610 (.Y(inst_cellmath__195[0]), .A0(N6554), .A1(N6052), .B0(N6252), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1611 (.Y(inst_cellmath__195[1]), .A0(N6554), .A1(N6204), .B0(N6403), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1612 (.Y(inst_cellmath__195[2]), .A0(N6554), .A1(N6362), .B0(N6555), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1613 (.Y(inst_cellmath__195[3]), .A0(N6554), .A1(N6508), .B0(N6008), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1614 (.Y(inst_cellmath__195[4]), .A0(N6554), .A1(N5953), .B0(N6162), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1615 (.Y(inst_cellmath__195[5]), .A0(N6554), .A1(N6114), .B0(N6317), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1616 (.Y(inst_cellmath__195[6]), .A0(N6554), .A1(N6269), .B0(N6462), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1617 (.Y(inst_cellmath__195[7]), .A0(N6554), .A1(N6416), .B0(N5909), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(inst_cellmath__195[8]), .A0(N6554), .A1(N6569), .B0(N6078), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1619 (.Y(inst_cellmath__195[9]), .A0(N6554), .A1(N6026), .B0(N6226), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1620 (.Y(inst_cellmath__195[10]), .A0(N6554), .A1(N6176), .B0(N6379), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1621 (.Y(inst_cellmath__195[11]), .A0(N6554), .A1(N6333), .B0(N6530), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1622 (.Y(inst_cellmath__195[12]), .A0(N6554), .A1(N6480), .B0(N5976), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1623 (.Y(inst_cellmath__195[13]), .A0(N6554), .A1(N5927), .B0(N6135), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1624 (.Y(inst_cellmath__195[14]), .A0(N6554), .A1(N6093), .B0(N6288), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1625 (.Y(inst_cellmath__195[15]), .A0(N6554), .A1(N6245), .B0(N6435), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1626 (.Y(inst_cellmath__195[16]), .A0(N6554), .A1(N6395), .B0(N5879), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1627 (.Y(inst_cellmath__195[17]), .A0(N6554), .A1(N6547), .B0(N6046), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1628 (.Y(inst_cellmath__195[18]), .A0(N6554), .A1(N5995), .B0(N6199), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1629 (.Y(inst_cellmath__195[19]), .A0(N6554), .A1(N6153), .B0(N6356), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1630 (.Y(inst_cellmath__195[20]), .A0(N6554), .A1(N6308), .B0(N6502), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1631 (.Y(inst_cellmath__195[21]), .A0(N6554), .A1(N6453), .B0(N5948), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1632 (.Y(inst_cellmath__195[22]), .A0(N6554), .A1(N5897), .B0(N6110), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1633 (.Y(inst_cellmath__195[23]), .A0(N6554), .A1(N6067), .B0(N6265), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1634 (.Y(inst_cellmath__195[24]), .A0(N6554), .A1(N6217), .B0(N6412), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1635 (.Y(inst_cellmath__195[25]), .A0(N6554), .A1(N6369), .B0(N6564), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1636 (.Y(inst_cellmath__195[26]), .A0(N6554), .A1(N6519), .B0(N6022), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1637 (.Y(inst_cellmath__195[27]), .A0(N6554), .A1(N5965), .B0(N6172), .B1(inst_cellmath__61[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1638 (.Y(inst_cellmath__195[28]), .A0(N6554), .A1(N6125), .B0(N5921), .B1(inst_cellmath__61[22]));
INVX1 inst_cellmath__198_0_I1640 (.Y(N7904), .A(inst_cellmath__61[1]));
INVXL inst_cellmath__198_0_I1641 (.Y(N7390), .A(inst_cellmath__61[2]));
INVXL inst_cellmath__198_0_I1642 (.Y(N7539), .A(inst_cellmath__61[3]));
INVXL inst_cellmath__198_0_I1643 (.Y(N7678), .A(inst_cellmath__61[4]));
INVXL inst_cellmath__198_0_I1644 (.Y(N7818), .A(inst_cellmath__61[5]));
INVXL inst_cellmath__198_0_I1645 (.Y(N7310), .A(inst_cellmath__61[6]));
INVXL inst_cellmath__198_0_I1646 (.Y(N7456), .A(inst_cellmath__61[7]));
INVXL inst_cellmath__198_0_I1647 (.Y(N7595), .A(inst_cellmath__61[8]));
INVXL inst_cellmath__198_0_I1648 (.Y(N7735), .A(inst_cellmath__61[9]));
INVXL inst_cellmath__198_0_I1649 (.Y(N7876), .A(inst_cellmath__61[10]));
INVXL inst_cellmath__198_0_I1650 (.Y(N7369), .A(inst_cellmath__61[11]));
INVXL inst_cellmath__198_0_I1651 (.Y(N7512), .A(inst_cellmath__61[12]));
INVXL inst_cellmath__198_0_I1652 (.Y(N7654), .A(inst_cellmath__61[13]));
INVXL inst_cellmath__198_0_I1653 (.Y(N7790), .A(inst_cellmath__61[14]));
INVXL inst_cellmath__198_0_I1654 (.Y(N7940), .A(inst_cellmath__61[15]));
INVXL inst_cellmath__198_0_I1655 (.Y(N7427), .A(inst_cellmath__115__W1[0]));
XOR2XL inst_cellmath__198_0_I8331 (.Y(N7570), .A(N684), .B(N5817));
NOR2XL inst_cellmath__198_0_I1660 (.Y(N7364), .A(N7570), .B(N7539));
NOR2XL inst_cellmath__198_0_I1661 (.Y(N7648), .A(N7570), .B(N7678));
NOR2XL inst_cellmath__198_0_I1662 (.Y(N7935), .A(N7570), .B(N7818));
NOR2XL inst_cellmath__198_0_I1663 (.Y(N7568), .A(N7570), .B(N7310));
NOR2XL inst_cellmath__198_0_I1664 (.Y(N7845), .A(N7570), .B(N7456));
NOR2XL inst_cellmath__198_0_I1665 (.Y(N7484), .A(N7570), .B(N7595));
NOR2XL inst_cellmath__198_0_I1666 (.Y(N7763), .A(N7570), .B(N7735));
NOR2XL inst_cellmath__198_0_I1667 (.Y(N7398), .A(N7570), .B(N7876));
NOR2XL inst_cellmath__198_0_I1668 (.Y(N7684), .A(N7570), .B(N7369));
NOR2XL inst_cellmath__198_0_I1669 (.Y(N7319), .A(N7570), .B(N7512));
NOR2XL inst_cellmath__198_0_I1670 (.Y(N7604), .A(N7570), .B(N7654));
NOR2XL inst_cellmath__198_0_I1671 (.Y(N7882), .A(N7570), .B(N7790));
NOR2XL inst_cellmath__198_0_I1672 (.Y(N7520), .A(N7570), .B(N7940));
OR2XL inst_cellmath__198_0_I1673 (.Y(N7565), .A(N7570), .B(N7427));
NOR2XL inst_cellmath__198_0_I1674 (.Y(N7469), .A(N7904), .B(N7390));
NOR2XL inst_cellmath__198_0_I1675 (.Y(N7749), .A(N7904), .B(N7539));
NOR2XL inst_cellmath__198_0_I1676 (.Y(N7383), .A(N7904), .B(N7678));
NOR2XL inst_cellmath__198_0_I1677 (.Y(N7670), .A(N7904), .B(N7818));
NOR2XL inst_cellmath__198_0_I1678 (.Y(N7304), .A(N7904), .B(N7310));
NOR2XL inst_cellmath__198_0_I1679 (.Y(N7588), .A(N7904), .B(N7456));
NOR2XL inst_cellmath__198_0_I1680 (.Y(N7867), .A(N7904), .B(N7595));
NOR2XL inst_cellmath__198_0_I1681 (.Y(N7505), .A(N7904), .B(N7735));
NOR2XL inst_cellmath__198_0_I1682 (.Y(N7782), .A(N7904), .B(N7876));
NOR2XL inst_cellmath__198_0_I1683 (.Y(N7419), .A(N7904), .B(N7369));
NOR2XL inst_cellmath__198_0_I1684 (.Y(N7705), .A(N7904), .B(N7512));
NOR2XL inst_cellmath__198_0_I1685 (.Y(N7339), .A(N7904), .B(N7654));
NOR2XL inst_cellmath__198_0_I1686 (.Y(N7625), .A(N7904), .B(N7790));
NOR2XL inst_cellmath__198_0_I1687 (.Y(N7908), .A(N7904), .B(N7940));
OR2XL inst_cellmath__198_0_I1688 (.Y(N7706), .A(N7904), .B(N7427));
INVXL inst_cellmath__198_0_I1689 (.Y(N7288), .A(N7390));
NOR2XL inst_cellmath__198_0_I1690 (.Y(N7851), .A(N7390), .B(N7539));
NOR2XL inst_cellmath__198_0_I1691 (.Y(N7490), .A(N7390), .B(N7678));
NOR2XL inst_cellmath__198_0_I1692 (.Y(N7768), .A(N7390), .B(N7818));
NOR2XL inst_cellmath__198_0_I1693 (.Y(N7404), .A(N7390), .B(N7310));
NOR2XL inst_cellmath__198_0_I1694 (.Y(N7690), .A(N7390), .B(N7456));
NOR2XL inst_cellmath__198_0_I1695 (.Y(N7324), .A(N7390), .B(N7595));
NOR2XL inst_cellmath__198_0_I1696 (.Y(N7610), .A(N7390), .B(N7735));
NOR2XL inst_cellmath__198_0_I1697 (.Y(N7889), .A(N7390), .B(N7876));
NOR2XL inst_cellmath__198_0_I1698 (.Y(N7525), .A(N7390), .B(N7369));
NOR2XL inst_cellmath__198_0_I1699 (.Y(N7805), .A(N7390), .B(N7512));
NOR2XL inst_cellmath__198_0_I1700 (.Y(N7442), .A(N7390), .B(N7654));
NOR2XL inst_cellmath__198_0_I1701 (.Y(N7725), .A(N7390), .B(N7790));
NOR2XL inst_cellmath__198_0_I1702 (.Y(N7358), .A(N7390), .B(N7940));
OR2XL inst_cellmath__198_0_I1703 (.Y(N7843), .A(N7390), .B(N7427));
INVXL inst_cellmath__198_0_I1704 (.Y(N7391), .A(N7539));
NOR2XL inst_cellmath__198_0_I1705 (.Y(N7311), .A(N7539), .B(N7678));
NOR2XL inst_cellmath__198_0_I1706 (.Y(N7596), .A(N7539), .B(N7818));
NOR2XL inst_cellmath__198_0_I1707 (.Y(N7875), .A(N7539), .B(N7310));
NOR2XL inst_cellmath__198_0_I1708 (.Y(N7513), .A(N7539), .B(N7456));
NOR2XL inst_cellmath__198_0_I1709 (.Y(N7791), .A(N7539), .B(N7595));
NOR2XL inst_cellmath__198_0_I1710 (.Y(N7426), .A(N7539), .B(N7735));
NOR2XL inst_cellmath__198_0_I1711 (.Y(N7712), .A(N7539), .B(N7876));
NOR2XL inst_cellmath__198_0_I1712 (.Y(N7346), .A(N7539), .B(N7369));
NOR2XL inst_cellmath__198_0_I1713 (.Y(N7631), .A(N7539), .B(N7512));
NOR2XL inst_cellmath__198_0_I1714 (.Y(N7915), .A(N7539), .B(N7654));
NOR2XL inst_cellmath__198_0_I1715 (.Y(N7549), .A(N7539), .B(N7790));
NOR2XL inst_cellmath__198_0_I1716 (.Y(N7826), .A(N7539), .B(N7940));
OR2XL inst_cellmath__198_0_I1717 (.Y(N7341), .A(N7539), .B(N7427));
INVXL inst_cellmath__198_0_I1718 (.Y(N7860), .A(N7678));
NOR2XL inst_cellmath__198_0_I1719 (.Y(N7776), .A(N7678), .B(N7818));
NOR2XL inst_cellmath__198_0_I1720 (.Y(N7413), .A(N7678), .B(N7310));
NOR2XL inst_cellmath__198_0_I1721 (.Y(N7698), .A(N7678), .B(N7456));
NOR2XL inst_cellmath__198_0_I1722 (.Y(N7332), .A(N7678), .B(N7595));
NOR2XL inst_cellmath__198_0_I1723 (.Y(N7619), .A(N7678), .B(N7735));
NOR2XL inst_cellmath__198_0_I1724 (.Y(N7899), .A(N7678), .B(N7876));
NOR2XL inst_cellmath__198_0_I1725 (.Y(N7534), .A(N7678), .B(N7369));
NOR2XL inst_cellmath__198_0_I1726 (.Y(N7813), .A(N7678), .B(N7512));
NOR2XL inst_cellmath__198_0_I1727 (.Y(N7451), .A(N7678), .B(N7654));
NOR2XL inst_cellmath__198_0_I1728 (.Y(N7730), .A(N7678), .B(N7790));
NOR2XL inst_cellmath__198_0_I1729 (.Y(N7365), .A(N7678), .B(N7940));
OR2XL inst_cellmath__198_0_I1730 (.Y(N7483), .A(N7678), .B(N7427));
INVXL inst_cellmath__198_0_I1731 (.Y(N7399), .A(N7818));
NOR2XL inst_cellmath__198_0_I1732 (.Y(N7320), .A(N7818), .B(N7310));
NOR2XL inst_cellmath__198_0_I1733 (.Y(N7606), .A(N7818), .B(N7456));
NOR2XL inst_cellmath__198_0_I1734 (.Y(N7885), .A(N7818), .B(N7595));
NOR2XL inst_cellmath__198_0_I1735 (.Y(N7522), .A(N7818), .B(N7735));
NOR2XL inst_cellmath__198_0_I1736 (.Y(N7800), .A(N7818), .B(N7876));
NOR2XL inst_cellmath__198_0_I1737 (.Y(N7437), .A(N7818), .B(N7369));
NOR2XL inst_cellmath__198_0_I1738 (.Y(N7720), .A(N7818), .B(N7512));
NOR2XL inst_cellmath__198_0_I1739 (.Y(N7354), .A(N7818), .B(N7654));
NOR2XL inst_cellmath__198_0_I1740 (.Y(N7639), .A(N7818), .B(N7790));
NOR2XL inst_cellmath__198_0_I1741 (.Y(N7924), .A(N7818), .B(N7940));
OR2XL inst_cellmath__198_0_I1742 (.Y(N7626), .A(N7818), .B(N7427));
INVXL inst_cellmath__198_0_I1743 (.Y(N7306), .A(N7310));
NOR2XL inst_cellmath__198_0_I1744 (.Y(N7869), .A(N7310), .B(N7456));
NOR2XL inst_cellmath__198_0_I1745 (.Y(N7507), .A(N7310), .B(N7595));
NOR2XL inst_cellmath__198_0_I1746 (.Y(N7785), .A(N7310), .B(N7735));
NOR2XL inst_cellmath__198_0_I1747 (.Y(N7421), .A(N7310), .B(N7876));
NOR2XL inst_cellmath__198_0_I1748 (.Y(N7707), .A(N7310), .B(N7369));
NOR2XL inst_cellmath__198_0_I1749 (.Y(N7342), .A(N7310), .B(N7512));
NOR2XL inst_cellmath__198_0_I1750 (.Y(N7628), .A(N7310), .B(N7654));
NOR2XL inst_cellmath__198_0_I1751 (.Y(N7911), .A(N7310), .B(N7790));
NOR2XL inst_cellmath__198_0_I1752 (.Y(N7545), .A(N7310), .B(N7940));
OR2XL inst_cellmath__198_0_I1753 (.Y(N7761), .A(N7310), .B(N7427));
INVXL inst_cellmath__198_0_I1754 (.Y(N7576), .A(N7456));
NOR2XL inst_cellmath__198_0_I1755 (.Y(N7494), .A(N7456), .B(N7595));
NOR2XL inst_cellmath__198_0_I1756 (.Y(N7770), .A(N7456), .B(N7735));
NOR2XL inst_cellmath__198_0_I1757 (.Y(N7407), .A(N7456), .B(N7876));
NOR2XL inst_cellmath__198_0_I1758 (.Y(N7694), .A(N7456), .B(N7369));
NOR2XL inst_cellmath__198_0_I1759 (.Y(N7325), .A(N7456), .B(N7512));
NOR2XL inst_cellmath__198_0_I1760 (.Y(N7613), .A(N7456), .B(N7654));
NOR2XL inst_cellmath__198_0_I1761 (.Y(N7893), .A(N7456), .B(N7790));
NOR2XL inst_cellmath__198_0_I1762 (.Y(N7527), .A(N7456), .B(N7940));
OR2XL inst_cellmath__198_0_I1763 (.Y(N7909), .A(N7456), .B(N7427));
INVXL inst_cellmath__198_0_I1764 (.Y(N7562), .A(N7595));
NOR2XL inst_cellmath__198_0_I1765 (.Y(N7480), .A(N7595), .B(N7735));
NOR2XL inst_cellmath__198_0_I1766 (.Y(N7759), .A(N7595), .B(N7876));
NOR2XL inst_cellmath__198_0_I1767 (.Y(N7394), .A(N7595), .B(N7369));
NOR2XL inst_cellmath__198_0_I1768 (.Y(N7680), .A(N7595), .B(N7512));
NOR2XL inst_cellmath__198_0_I1769 (.Y(N7314), .A(N7595), .B(N7654));
NOR2XL inst_cellmath__198_0_I1770 (.Y(N7599), .A(N7595), .B(N7790));
NOR2XL inst_cellmath__198_0_I1771 (.Y(N7878), .A(N7595), .B(N7940));
OR2XL inst_cellmath__198_0_I1772 (.Y(N7395), .A(N7595), .B(N7427));
INVXL inst_cellmath__198_0_I1773 (.Y(N7918), .A(N7735));
NOR2XL inst_cellmath__198_0_I1774 (.Y(N7828), .A(N7735), .B(N7876));
NOR2XL inst_cellmath__198_0_I1775 (.Y(N7465), .A(N7735), .B(N7369));
NOR2XL inst_cellmath__198_0_I1776 (.Y(N7745), .A(N7735), .B(N7512));
NOR2XL inst_cellmath__198_0_I1777 (.Y(N7379), .A(N7735), .B(N7654));
NOR2XL inst_cellmath__198_0_I1778 (.Y(N7665), .A(N7735), .B(N7790));
NOR2XL inst_cellmath__198_0_I1779 (.Y(N7300), .A(N7735), .B(N7940));
OR2XL inst_cellmath__198_0_I1780 (.Y(N7543), .A(N7735), .B(N7427));
INVXL inst_cellmath__198_0_I1781 (.Y(N7336), .A(N7876));
NOR2XL inst_cellmath__198_0_I1782 (.Y(N7903), .A(N7876), .B(N7369));
NOR2XL inst_cellmath__198_0_I1783 (.Y(N7538), .A(N7876), .B(N7512));
NOR2XL inst_cellmath__198_0_I1784 (.Y(N7817), .A(N7876), .B(N7654));
NOR2XL inst_cellmath__198_0_I1785 (.Y(N7455), .A(N7876), .B(N7790));
NOR2XL inst_cellmath__198_0_I1786 (.Y(N7734), .A(N7876), .B(N7940));
OR2XL inst_cellmath__198_0_I1787 (.Y(N7682), .A(N7876), .B(N7427));
INVXL inst_cellmath__198_0_I1788 (.Y(N7765), .A(N7369));
NOR2XL inst_cellmath__198_0_I1789 (.Y(N7687), .A(N7369), .B(N7512));
NOR2XL inst_cellmath__198_0_I1790 (.Y(N7322), .A(N7369), .B(N7654));
NOR2XL inst_cellmath__198_0_I1791 (.Y(N7608), .A(N7369), .B(N7790));
NOR2XL inst_cellmath__198_0_I1792 (.Y(N7887), .A(N7369), .B(N7940));
OR2XL inst_cellmath__198_0_I1793 (.Y(N7822), .A(N7369), .B(N7427));
INVXL inst_cellmath__198_0_I1794 (.Y(N7926), .A(N7512));
NOR2XL inst_cellmath__198_0_I1795 (.Y(N7837), .A(N7512), .B(N7654));
NOR2XL inst_cellmath__198_0_I1796 (.Y(N7473), .A(N7512), .B(N7790));
NOR2XL inst_cellmath__198_0_I1797 (.Y(N7753), .A(N7512), .B(N7940));
OR2XL inst_cellmath__198_0_I1798 (.Y(N7316), .A(N7512), .B(N7427));
INVXL inst_cellmath__198_0_I1799 (.Y(N7787), .A(N7654));
NOR2XL inst_cellmath__198_0_I1800 (.Y(N7709), .A(N7654), .B(N7790));
NOR2XL inst_cellmath__198_0_I1801 (.Y(N7344), .A(N7654), .B(N7940));
OR2XL inst_cellmath__198_0_I1802 (.Y(N7459), .A(N7654), .B(N7427));
INVXL inst_cellmath__198_0_I1803 (.Y(N7375), .A(N7790));
NOR2XL inst_cellmath__198_0_I1804 (.Y(N7293), .A(N7790), .B(N7940));
OR2XL inst_cellmath__198_0_I1805 (.Y(N7601), .A(N7790), .B(N7427));
INVXL inst_cellmath__198_0_I1806 (.Y(N7328), .A(N7940));
ADDHX1 inst_cellmath__198_0_I1807 (.CO(N7880), .S(N7739), .A(N7684), .B(N7320));
ADDHX1 inst_cellmath__198_0_I1808 (.CO(N7517), .S(N7372), .A(N7419), .B(N7606));
ADDFX1 inst_cellmath__198_0_I1809 (.CO(N7795), .S(N7657), .A(N7604), .B(N7576), .CI(N7885));
ADDHX1 inst_cellmath__198_0_I1810 (.CO(N7431), .S(N7290), .A(N7712), .B(N7705));
ADDFX1 inst_cellmath__198_0_I1811 (.CO(N7716), .S(N7574), .A(N7522), .B(N7339), .CI(N7346));
ADDHX1 inst_cellmath__198_0_I1812 (.CO(N7349), .S(N7852), .A(N7882), .B(N7507));
ADDFX1 inst_cellmath__198_0_I1813 (.CO(N7635), .S(N7492), .A(N7562), .B(N7520), .CI(N7494));
ADDFX1 inst_cellmath__198_0_I1814 (.CO(N7920), .S(N7769), .A(N7631), .B(N7800), .CI(N7625));
ADDHX1 inst_cellmath__198_0_I1815 (.CO(N7552), .S(N7405), .A(N7785), .B(N7534));
XNOR2X1 inst_cellmath__198_0_I1816 (.Y(N7692), .A(N7908), .B(N7770));
OR2XL inst_cellmath__198_0_I1817 (.Y(N7830), .A(N7908), .B(N7770));
ADDFX1 inst_cellmath__198_0_I1818 (.CO(N7746), .S(N7611), .A(N7915), .B(N7437), .CI(N7565));
ADDFX1 inst_cellmath__198_0_I1819 (.CO(N7380), .S(N7891), .A(N7813), .B(N7421), .CI(N7725));
ADDFX1 inst_cellmath__198_0_I1820 (.CO(N7667), .S(N7526), .A(N7706), .B(N7918), .CI(N7407));
ADDFX1 inst_cellmath__198_0_I1821 (.CO(N7301), .S(N7806), .A(N7549), .B(N7720), .CI(N7480));
ADDFX1 inst_cellmath__198_0_I1822 (.CO(N7586), .S(N7444), .A(N7451), .B(N7707), .CI(N7358));
ADDFX1 inst_cellmath__198_0_I1823 (.CO(N7865), .S(N7726), .A(N7354), .B(N7694), .CI(N7826));
ADDFX1 inst_cellmath__198_0_I1824 (.CO(N7503), .S(N7359), .A(N7342), .B(N7759), .CI(N7730));
ADDFX1 inst_cellmath__198_0_I1825 (.CO(N7780), .S(N7643), .A(N7341), .B(N7336), .CI(N7828));
ADDFX1 inst_cellmath__198_0_I1826 (.CO(N7417), .S(N7931), .A(N7639), .B(N7325), .CI(N7394));
ADDFX1 inst_cellmath__198_0_I1827 (.CO(N7702), .S(N7560), .A(N7613), .B(N7465), .CI(N7924));
ADDFX1 inst_cellmath__198_0_I1828 (.CO(N7337), .S(N7841), .A(N7626), .B(N7765), .CI(N7745));
ADDHX1 inst_cellmath__198_0_I1829 (.CO(N7623), .S(N7479), .A(N7845), .B(N7311));
ADDHX1 inst_cellmath__198_0_I1830 (.CO(N7906), .S(N7757), .A(N7588), .B(N7596));
ADDFX1 inst_cellmath__198_0_I1831 (.CO(N7540), .S(N7392), .A(N7763), .B(N7399), .CI(N7875));
ADDHX1 inst_cellmath__198_0_I1832 (.CO(N7819), .S(N7679), .A(N7867), .B(N7776));
ADDFX1 inst_cellmath__198_0_I1833 (.CO(N7457), .S(N7312), .A(N7513), .B(N7505), .CI(N7398));
ADDHX1 inst_cellmath__198_0_I1834 (.CO(N7736), .S(N7597), .A(N7413), .B(N7324));
ADDFX1 inst_cellmath__198_0_I1835 (.CO(N7370), .S(N7877), .A(N7791), .B(N7306), .CI(N7782));
ADDFX1 inst_cellmath__198_0_I1836 (.CO(N7655), .S(N7514), .A(N7610), .B(N7698), .CI(N7739));
ADDFX1 inst_cellmath__198_0_I1837 (.CO(N7286), .S(N7792), .A(N7319), .B(N7426), .CI(N7332));
ADDFX1 inst_cellmath__198_0_I1838 (.CO(N7572), .S(N7428), .A(N7880), .B(N7889), .CI(N7372));
ADDFX1 inst_cellmath__198_0_I1839 (.CO(N7849), .S(N7713), .A(N7619), .B(N7869), .CI(N7525));
ADDFX1 inst_cellmath__198_0_I1840 (.CO(N7488), .S(N7347), .A(N7290), .B(N7517), .CI(N7657));
ADDFX1 inst_cellmath__198_0_I1841 (.CO(N7766), .S(N7633), .A(N7805), .B(N7899), .CI(N7431));
ADDFX1 inst_cellmath__198_0_I1842 (.CO(N7402), .S(N7916), .A(N7852), .B(N7795), .CI(N7574));
ADDFX1 inst_cellmath__198_0_I1843 (.CO(N7688), .S(N7550), .A(N7349), .B(N7442), .CI(N7716));
ADDFX1 inst_cellmath__198_0_I1844 (.CO(N7323), .S(N7827), .A(N7492), .B(N7405), .CI(N7769));
ADDFX1 inst_cellmath__198_0_I1845 (.CO(N7609), .S(N7464), .A(N7692), .B(N7552), .CI(N7635));
ADDFX1 inst_cellmath__198_0_I1846 (.CO(N7888), .S(N7744), .A(N7611), .B(N7920), .CI(N7891));
ADDFX1 inst_cellmath__198_0_I1847 (.CO(N7524), .S(N7378), .A(N7746), .B(N7830), .CI(N7380));
ADDFX1 inst_cellmath__198_0_I1848 (.CO(N7804), .S(N7663), .A(N7806), .B(N7526), .CI(N7444));
ADDFX1 inst_cellmath__198_0_I1849 (.CO(N7440), .S(N7297), .A(N7667), .B(N7843), .CI(N7301));
ADDFX1 inst_cellmath__198_0_I1850 (.CO(N7723), .S(N7582), .A(N7726), .B(N7586), .CI(N7359));
ADDFX1 inst_cellmath__198_0_I1851 (.CO(N7356), .S(N7861), .A(N7365), .B(N7628), .CI(N7865));
ADDFX1 inst_cellmath__198_0_I1852 (.CO(N7641), .S(N7500), .A(N7643), .B(N7503), .CI(N7931));
ADDFX1 inst_cellmath__198_0_I1853 (.CO(N7927), .S(N7777), .A(N7911), .B(N7680), .CI(N7483));
ADDFX1 inst_cellmath__198_0_I1854 (.CO(N7557), .S(N7414), .A(N7417), .B(N7780), .CI(N7560));
ADDFX1 inst_cellmath__198_0_I1855 (.CO(N7838), .S(N7699), .A(N7903), .B(N7893), .CI(N7314));
ADDFX1 inst_cellmath__198_0_I1856 (.CO(N7476), .S(N7333), .A(N7702), .B(N7545), .CI(N7841));
ADDFX1 inst_cellmath__198_0_I1857 (.CO(N7754), .S(N7620), .A(N7527), .B(N7379), .CI(N7538));
ADDFX1 inst_cellmath__198_0_I1858 (.CO(N7388), .S(N7900), .A(N7761), .B(N7599), .CI(N7337));
ADDFX1 inst_cellmath__198_0_I1859 (.CO(N7676), .S(N7535), .A(N7909), .B(N7926), .CI(N7687));
ADDFX1 inst_cellmath__198_0_I1860 (.CO(N7308), .S(N7814), .A(N7817), .B(N7665), .CI(N7878));
ADDFX1 inst_cellmath__198_0_I1861 (.CO(N7592), .S(N7452), .A(N7300), .B(N7322), .CI(N7455));
ADDFX1 inst_cellmath__198_0_I1862 (.CO(N7872), .S(N7731), .A(N7543), .B(N7787), .CI(N7608));
ADDHX1 inst_cellmath__198_0_I1863 (.CO(N7509), .S(N7366), .A(N7935), .B(N7391));
ADDHX1 inst_cellmath__198_0_I1864 (.CO(N7788), .S(N7650), .A(N7670), .B(N7568));
ADDFX1 inst_cellmath__198_0_I1865 (.CO(N7424), .S(N7938), .A(N7860), .B(N7304), .CI(N7768));
ADDFX1 inst_cellmath__198_0_I1866 (.CO(N7710), .S(N7569), .A(N7404), .B(N7484), .CI(N7623));
ADDFX1 inst_cellmath__198_0_I1867 (.CO(N7345), .S(N7847), .A(N7906), .B(N7690), .CI(N7679));
ADDFX1 inst_cellmath__198_0_I1868 (.CO(N7630), .S(N7486), .A(N7540), .B(N7819), .CI(N7597));
ADDFX1 inst_cellmath__198_0_I1869 (.CO(N7914), .S(N7764), .A(N7457), .B(N7736), .CI(N7877));
ADDFX1 inst_cellmath__198_0_I1870 (.CO(N7547), .S(N7400), .A(N7792), .B(N7370), .CI(N7655));
ADDFX1 inst_cellmath__198_0_I1871 (.CO(N7825), .S(N7686), .A(N7572), .B(N7286), .CI(N7713));
ADDFX1 inst_cellmath__198_0_I1872 (.CO(N7463), .S(N7321), .A(N7633), .B(N7849), .CI(N7488));
ADDFX1 inst_cellmath__198_0_I1873 (.CO(N7742), .S(N7607), .A(N7402), .B(N7766), .CI(N7550));
ADDFX1 inst_cellmath__198_0_I1874 (.CO(N7377), .S(N7886), .A(N7464), .B(N7688), .CI(N7323));
ADDFX1 inst_cellmath__198_0_I1875 (.CO(N7661), .S(N7523), .A(N7378), .B(N7609), .CI(N7888));
ADDFX1 inst_cellmath__198_0_I1876 (.CO(N7296), .S(N7801), .A(N7297), .B(N7524), .CI(N7804));
ADDFX1 inst_cellmath__198_0_I1877 (.CO(N7581), .S(N7438), .A(N7861), .B(N7440), .CI(N7723));
ADDFX1 inst_cellmath__198_0_I1878 (.CO(N7859), .S(N7722), .A(N7777), .B(N7356), .CI(N7641));
ADDFX1 inst_cellmath__198_0_I1879 (.CO(N7499), .S(N7355), .A(N7699), .B(N7927), .CI(N7557));
ADDFX1 inst_cellmath__198_0_I1880 (.CO(N7775), .S(N7640), .A(N7620), .B(N7838), .CI(N7476));
ADDFX1 inst_cellmath__198_0_I1881 (.CO(N7411), .S(N7925), .A(N7535), .B(N7754), .CI(N7814));
ADDFX1 inst_cellmath__198_0_I1882 (.CO(N7697), .S(N7556), .A(N7676), .B(N7395), .CI(N7308));
ADDFX1 inst_cellmath__198_0_I1883 (.CO(N7330), .S(N7835), .A(N7734), .B(N7837), .CI(N7592));
ADDFX1 inst_cellmath__198_0_I1884 (.CO(N7616), .S(N7471), .A(N7473), .B(N7887), .CI(N7682));
ADDFX1 inst_cellmath__198_0_I1885 (.CO(N7896), .S(N7751), .A(N7822), .B(N7375), .CI(N7709));
ADDHX1 inst_cellmath__198_0_I1886 (.CO(N7532), .S(N7386), .A(N7364), .B(N7469));
ADDHX1 inst_cellmath__198_0_I1887 (.CO(N7811), .S(N7672), .A(N7749), .B(N7648));
ADDFX1 inst_cellmath__198_0_I1888 (.CO(N7448), .S(N7307), .A(N7851), .B(N7383), .CI(N7366));
ADDFX1 inst_cellmath__198_0_I1889 (.CO(N7729), .S(N7591), .A(N7509), .B(N7490), .CI(N7650));
ADDFX1 inst_cellmath__198_0_I1890 (.CO(N7363), .S(N7870), .A(N7479), .B(N7788), .CI(N7938));
ADDFX1 inst_cellmath__198_0_I1891 (.CO(N7647), .S(N7508), .A(N7424), .B(N7757), .CI(N7569));
ADDFX1 inst_cellmath__198_0_I1892 (.CO(N7936), .S(N7786), .A(N7392), .B(N7710), .CI(N7847));
ADDFX1 inst_cellmath__198_0_I1893 (.CO(N7567), .S(N7422), .A(N7345), .B(N7312), .CI(N7486));
ADDFX1 inst_cellmath__198_0_I1894 (.CO(N7844), .S(N7708), .A(N7514), .B(N7630), .CI(N7764));
ADDFX1 inst_cellmath__198_0_I1895 (.CO(N7485), .S(N7343), .A(N7914), .B(N7428), .CI(N7400));
ADDFX1 inst_cellmath__198_0_I1896 (.CO(N7762), .S(N7629), .A(N7347), .B(N7547), .CI(N7686));
ADDFX1 inst_cellmath__198_0_I1897 (.CO(N7397), .S(N7912), .A(N7916), .B(N7825), .CI(N7321));
ADDFX1 inst_cellmath__198_0_I1898 (.CO(N7685), .S(N7546), .A(N7463), .B(N7827), .CI(N7607));
ADDFX1 inst_cellmath__198_0_I1899 (.CO(N7318), .S(N7824), .A(N7742), .B(N7744), .CI(N7886));
ADDFX1 inst_cellmath__198_0_I1900 (.CO(N7603), .S(N7462), .A(N7377), .B(N7663), .CI(N7523));
ADDFX1 inst_cellmath__198_0_I1901 (.CO(N7883), .S(N7741), .A(N7661), .B(N7582), .CI(N7801));
ADDFX1 inst_cellmath__198_0_I1902 (.CO(N7519), .S(N7374), .A(N7296), .B(N7500), .CI(N7438));
ADDFX1 inst_cellmath__198_0_I1903 (.CO(N7797), .S(N7659), .A(N7581), .B(N7414), .CI(N7722));
ADDFX1 inst_cellmath__198_0_I1904 (.CO(N7434), .S(N7292), .A(N7859), .B(N7333), .CI(N7355));
ADDFX1 inst_cellmath__198_0_I1905 (.CO(N7718), .S(N7577), .A(N7499), .B(N7900), .CI(N7640));
ADDFX1 inst_cellmath__198_0_I1906 (.CO(N7351), .S(N7854), .A(N7925), .B(N7388), .CI(N7775));
ADDFX1 inst_cellmath__198_0_I1907 (.CO(N7637), .S(N7495), .A(N7556), .B(N7452), .CI(N7411));
ADDFX1 inst_cellmath__198_0_I1908 (.CO(N7922), .S(N7772), .A(N7697), .B(N7731), .CI(N7835));
ADDFX1 inst_cellmath__198_0_I1909 (.CO(N7554), .S(N7408), .A(N7471), .B(N7872), .CI(N7330));
ADDFX1 inst_cellmath__198_0_I1910 (.CO(N7832), .S(N7695), .A(N7616), .B(N7753), .CI(N7751));
ADDFX1 inst_cellmath__198_0_I1911 (.CO(N7468), .S(N7327), .A(N7316), .B(N7344), .CI(N7896));
ADDFX1 inst_cellmath__198_0_I1912 (.CO(N7748), .S(N7614), .A(N7459), .B(N7328), .CI(N7293));
AND2XL inst_cellmath__198_0_I1915 (.Y(N7669), .A(N7288), .B(N7386));
NOR2XL inst_cellmath__198_0_I1916 (.Y(N7808), .A(N7532), .B(N7672));
NAND2XL inst_cellmath__198_0_I1917 (.Y(N7303), .A(N7532), .B(N7672));
AND2XL inst_cellmath__198_0_I1919 (.Y(N7587), .A(N7811), .B(N7307));
NOR2XL inst_cellmath__198_0_I1920 (.Y(N7727), .A(N7448), .B(N7591));
NAND2XL inst_cellmath__198_0_I1921 (.Y(N7866), .A(N7448), .B(N7591));
AND2XL inst_cellmath__198_0_I1923 (.Y(N7504), .A(N7729), .B(N7870));
NOR2XL inst_cellmath__198_0_I1924 (.Y(N7645), .A(N7363), .B(N7508));
NAND2XL inst_cellmath__198_0_I1925 (.Y(N7781), .A(N7363), .B(N7508));
NOR2XL inst_cellmath__198_0_I1926 (.Y(N7933), .A(N7647), .B(N7786));
NOR2XL inst_cellmath__198_0_I1928 (.Y(N7563), .A(N7936), .B(N7422));
NAND2XL inst_cellmath__198_0_I1929 (.Y(N7704), .A(N7936), .B(N7422));
NOR3XL inst_cellmath__198_0_I8376 (.Y(N7482), .A(N7570), .B(N7904), .C(N7390));
OAI22XL inst_cellmath__198_0_I8334 (.Y(N7600), .A0(N7669), .A1(N7482), .B0(N7288), .B1(N7386));
AOI21XL inst_cellmath__198_0_I1934 (.Y(N7430), .A0(N7303), .A1(N7600), .B0(N7808));
OAI22XL inst_cellmath__198_0_I8335 (.Y(N7829), .A0(N7587), .A1(N7430), .B0(N7811), .B1(N7307));
AOI21XL inst_cellmath__198_0_I1938 (.Y(N7585), .A0(N7866), .A1(N7829), .B0(N7727));
OAI22XL inst_cellmath__198_0_I8336 (.Y(N7905), .A0(N7504), .A1(N7585), .B0(N7729), .B1(N7870));
AOI21XL inst_cellmath__198_0_I1942 (.Y(N7571), .A0(N7781), .A1(N7905), .B0(N7645));
AOI21XL inst_cellmath__198_0_I1945 (.Y(N7487), .A0(N7704), .A1(N7933), .B0(N7563));
OAI2BB1X1 inst_cellmath__198_0_I8337 (.Y(N7632), .A0N(N7647), .A1N(N7786), .B0(N7704));
OAI21XL inst_cellmath__198_0_I1948 (.Y(N7605), .A0(N7632), .A1(N7571), .B0(N7487));
NOR2XL inst_cellmath__198_0_I1967 (.Y(N7884), .A(N7567), .B(N7708));
NAND2XL inst_cellmath__198_0_I1968 (.Y(N7376), .A(N7567), .B(N7708));
NOR2XL inst_cellmath__198_0_I1969 (.Y(N7521), .A(N7844), .B(N7343));
NAND2XL inst_cellmath__198_0_I1970 (.Y(N7660), .A(N7844), .B(N7343));
NOR2XL inst_cellmath__198_0_I1971 (.Y(N7799), .A(N7485), .B(N7629));
NAND2XL inst_cellmath__198_0_I1972 (.Y(N7294), .A(N7485), .B(N7629));
NOR2XL inst_cellmath__198_0_I1973 (.Y(N7436), .A(N7762), .B(N7912));
NAND2XL inst_cellmath__198_0_I1974 (.Y(N7580), .A(N7762), .B(N7912));
NOR2XL inst_cellmath__198_0_I1975 (.Y(N7719), .A(N7397), .B(N7546));
NAND2XL inst_cellmath__198_0_I1976 (.Y(N7858), .A(N7397), .B(N7546));
NOR2XL inst_cellmath__198_0_I1977 (.Y(N7353), .A(N7685), .B(N7824));
NAND2XL inst_cellmath__198_0_I1978 (.Y(N7497), .A(N7685), .B(N7824));
NOR2XL inst_cellmath__198_0_I1979 (.Y(N7638), .A(N7318), .B(N7462));
NAND2XL inst_cellmath__198_0_I1980 (.Y(N7774), .A(N7318), .B(N7462));
NOR2XL inst_cellmath__198_0_I1981 (.Y(N7923), .A(N7603), .B(N7741));
NAND2XL inst_cellmath__198_0_I1982 (.Y(N7410), .A(N7603), .B(N7741));
NOR2XL inst_cellmath__198_0_I1983 (.Y(N7555), .A(N7883), .B(N7374));
NAND2XL inst_cellmath__198_0_I1984 (.Y(N7696), .A(N7883), .B(N7374));
NOR2XL inst_cellmath__198_0_I1985 (.Y(N7833), .A(N7519), .B(N7659));
NAND2XL inst_cellmath__198_0_I1986 (.Y(N7329), .A(N7519), .B(N7659));
NOR2XL inst_cellmath__198_0_I1987 (.Y(N7470), .A(N7797), .B(N7292));
NAND2XL inst_cellmath__198_0_I1988 (.Y(N7615), .A(N7797), .B(N7292));
NOR2XL inst_cellmath__198_0_I1989 (.Y(N7750), .A(N7434), .B(N7577));
NAND2XL inst_cellmath__198_0_I1990 (.Y(N7895), .A(N7434), .B(N7577));
NOR2XL inst_cellmath__198_0_I1991 (.Y(N7385), .A(N7854), .B(N7718));
NAND2XL inst_cellmath__198_0_I1992 (.Y(N7531), .A(N7854), .B(N7718));
NOR2XL inst_cellmath__198_0_I1993 (.Y(N7671), .A(N7495), .B(N7351));
NAND2XL inst_cellmath__198_0_I1994 (.Y(N7810), .A(N7495), .B(N7351));
NOR2XL inst_cellmath__198_0_I1995 (.Y(N7305), .A(N7637), .B(N7772));
NAND2XL inst_cellmath__198_0_I1996 (.Y(N7447), .A(N7637), .B(N7772));
NOR2XL inst_cellmath__198_0_I1997 (.Y(N7590), .A(N7408), .B(N7922));
NAND2XL inst_cellmath__198_0_I1998 (.Y(N7728), .A(N7408), .B(N7922));
NOR2XL inst_cellmath__198_0_I1999 (.Y(N7868), .A(N7554), .B(N7695));
NAND2XL inst_cellmath__198_0_I2000 (.Y(N7362), .A(N7554), .B(N7695));
NOR2XL inst_cellmath__198_0_I2001 (.Y(N7506), .A(N7327), .B(N7832));
NAND2XL inst_cellmath__198_0_I2002 (.Y(N7646), .A(N7327), .B(N7832));
NOR2XL inst_cellmath__198_0_I2003 (.Y(N7784), .A(N7614), .B(N7468));
NAND2XL inst_cellmath__198_0_I2004 (.Y(N7934), .A(N7614), .B(N7468));
NOR2XL inst_cellmath__198_0_I2005 (.Y(N7420), .A(N7601), .B(N7748));
NAND2XL inst_cellmath__198_0_I2006 (.Y(N7566), .A(N7601), .B(N7748));
AO21XL inst_cellmath__198_0_I2007 (.Y(N7627), .A0(N7376), .A1(N7605), .B0(N7884));
AO21XL inst_cellmath__198_0_I2008 (.Y(N7910), .A0(N7660), .A1(N7884), .B0(N7521));
AND2XL inst_cellmath__198_0_I2009 (.Y(N7396), .A(N7660), .B(N7376));
AO21XL inst_cellmath__198_0_I2010 (.Y(N7544), .A0(N7294), .A1(N7521), .B0(N7799));
AND2XL inst_cellmath__198_0_I2011 (.Y(N7683), .A(N7294), .B(N7660));
AO21XL inst_cellmath__198_0_I2012 (.Y(N7823), .A0(N7580), .A1(N7799), .B0(N7436));
AND2XL inst_cellmath__198_0_I2013 (.Y(N7317), .A(N7580), .B(N7294));
AO21XL inst_cellmath__198_0_I2014 (.Y(N7460), .A0(N7858), .A1(N7436), .B0(N7719));
AND2XL inst_cellmath__198_0_I2015 (.Y(N7602), .A(N7858), .B(N7580));
AO21XL inst_cellmath__198_0_I2016 (.Y(N7740), .A0(N7497), .A1(N7719), .B0(N7353));
AND2XL inst_cellmath__198_0_I2017 (.Y(N7881), .A(N7497), .B(N7858));
AO21XL inst_cellmath__198_0_I2018 (.Y(N7373), .A0(N7774), .A1(N7353), .B0(N7638));
AND2XL inst_cellmath__198_0_I2019 (.Y(N7518), .A(N7774), .B(N7497));
AO21XL inst_cellmath__198_0_I2020 (.Y(N7658), .A0(N7410), .A1(N7638), .B0(N7923));
AND2XL inst_cellmath__198_0_I2021 (.Y(N7796), .A(N7410), .B(N7774));
AO21XL inst_cellmath__198_0_I2022 (.Y(N7291), .A0(N7696), .A1(N7923), .B0(N7555));
AND2XL inst_cellmath__198_0_I2023 (.Y(N7432), .A(N7696), .B(N7410));
AO21XL inst_cellmath__198_0_I2024 (.Y(N7575), .A0(N7329), .A1(N7555), .B0(N7833));
AND2XL inst_cellmath__198_0_I2025 (.Y(N7717), .A(N7329), .B(N7696));
AO21XL inst_cellmath__198_0_I2026 (.Y(N7853), .A0(N7615), .A1(N7833), .B0(N7470));
AND2XL inst_cellmath__198_0_I2027 (.Y(N7350), .A(N7615), .B(N7329));
AO21XL inst_cellmath__198_0_I2028 (.Y(N7493), .A0(N7895), .A1(N7470), .B0(N7750));
AND2XL inst_cellmath__198_0_I2029 (.Y(N7636), .A(N7895), .B(N7615));
AO21XL inst_cellmath__198_0_I2030 (.Y(N7771), .A0(N7531), .A1(N7750), .B0(N7385));
AND2XL inst_cellmath__198_0_I2031 (.Y(N7921), .A(N7531), .B(N7895));
AO21XL inst_cellmath__198_0_I2032 (.Y(N7406), .A0(N7810), .A1(N7385), .B0(N7671));
AND2XL inst_cellmath__198_0_I2033 (.Y(N7553), .A(N7810), .B(N7531));
AO21XL inst_cellmath__198_0_I2034 (.Y(N7693), .A0(N7447), .A1(N7671), .B0(N7305));
AND2XL inst_cellmath__198_0_I2035 (.Y(N7831), .A(N7447), .B(N7810));
AO21XL inst_cellmath__198_0_I2036 (.Y(N7326), .A0(N7728), .A1(N7305), .B0(N7590));
AND2XL inst_cellmath__198_0_I2037 (.Y(N7467), .A(N7728), .B(N7447));
AO21XL inst_cellmath__198_0_I2038 (.Y(N7612), .A0(N7362), .A1(N7590), .B0(N7868));
AND2XL inst_cellmath__198_0_I2039 (.Y(N7747), .A(N7362), .B(N7728));
AO21XL inst_cellmath__198_0_I2040 (.Y(N7892), .A0(N7646), .A1(N7868), .B0(N7506));
AND2XL inst_cellmath__198_0_I2041 (.Y(N7381), .A(N7646), .B(N7362));
AO21XL inst_cellmath__198_0_I2042 (.Y(N7528), .A0(N7934), .A1(N7506), .B0(N7784));
AND2XL inst_cellmath__198_0_I2043 (.Y(N7668), .A(N7934), .B(N7646));
AO21XL inst_cellmath__198_0_I2044 (.Y(N7807), .A0(N7566), .A1(N7784), .B0(N7420));
AND2XL inst_cellmath__198_0_I2045 (.Y(N7302), .A(N7566), .B(N7934));
AO21XL inst_cellmath__198_0_I2046 (.Y(N7644), .A0(N7605), .A1(N7396), .B0(N7910));
AO21XL inst_cellmath__198_0_I2047 (.Y(N7932), .A0(N7683), .A1(N7627), .B0(N7544));
AO21XL inst_cellmath__198_0_I2048 (.Y(N7561), .A0(N7317), .A1(N7910), .B0(N7823));
AND2XL inst_cellmath__198_0_I2049 (.Y(N7703), .A(N7317), .B(N7396));
AO21XL inst_cellmath__198_0_I2050 (.Y(N7842), .A0(N7602), .A1(N7544), .B0(N7460));
AND2XL inst_cellmath__198_0_I2051 (.Y(N7338), .A(N7602), .B(N7683));
AO21XL inst_cellmath__198_0_I2052 (.Y(N7481), .A0(N7881), .A1(N7823), .B0(N7740));
AND2XL inst_cellmath__198_0_I2053 (.Y(N7624), .A(N7881), .B(N7317));
AO21XL inst_cellmath__198_0_I2054 (.Y(N7758), .A0(N7518), .A1(N7460), .B0(N7373));
AND2XL inst_cellmath__198_0_I2055 (.Y(N7907), .A(N7518), .B(N7602));
AO21XL inst_cellmath__198_0_I2056 (.Y(N7393), .A0(N7796), .A1(N7740), .B0(N7658));
AND2XL inst_cellmath__198_0_I2057 (.Y(N7541), .A(N7796), .B(N7881));
AO21XL inst_cellmath__198_0_I2058 (.Y(N7681), .A0(N7432), .A1(N7373), .B0(N7291));
AND2XL inst_cellmath__198_0_I2059 (.Y(N7820), .A(N7432), .B(N7518));
AO21XL inst_cellmath__198_0_I2060 (.Y(N7313), .A0(N7717), .A1(N7658), .B0(N7575));
AND2XL inst_cellmath__198_0_I2061 (.Y(N7458), .A(N7717), .B(N7796));
AO21XL inst_cellmath__198_0_I2062 (.Y(N7598), .A0(N7350), .A1(N7291), .B0(N7853));
AND2XL inst_cellmath__198_0_I2063 (.Y(N7737), .A(N7350), .B(N7432));
AO21XL inst_cellmath__198_0_I2064 (.Y(N7879), .A0(N7636), .A1(N7575), .B0(N7493));
AND2XL inst_cellmath__198_0_I2065 (.Y(N7371), .A(N7636), .B(N7717));
AO21XL inst_cellmath__198_0_I2066 (.Y(N7515), .A0(N7921), .A1(N7853), .B0(N7771));
AND2XL inst_cellmath__198_0_I2067 (.Y(N7656), .A(N7921), .B(N7350));
AO21XL inst_cellmath__198_0_I2068 (.Y(N7793), .A0(N7553), .A1(N7493), .B0(N7406));
AND2XL inst_cellmath__198_0_I2069 (.Y(N7287), .A(N7553), .B(N7636));
AO21XL inst_cellmath__198_0_I2070 (.Y(N7429), .A0(N7831), .A1(N7771), .B0(N7693));
AND2XL inst_cellmath__198_0_I2071 (.Y(N7573), .A(N7831), .B(N7921));
AO21XL inst_cellmath__198_0_I2072 (.Y(N7714), .A0(N7467), .A1(N7406), .B0(N7326));
AND2XL inst_cellmath__198_0_I2073 (.Y(N7850), .A(N7467), .B(N7553));
AO21XL inst_cellmath__198_0_I2074 (.Y(N7348), .A0(N7747), .A1(N7693), .B0(N7612));
AND2XL inst_cellmath__198_0_I2075 (.Y(N7489), .A(N7747), .B(N7831));
AO21XL inst_cellmath__198_0_I2076 (.Y(N7634), .A0(N7381), .A1(N7326), .B0(N7892));
AND2XL inst_cellmath__198_0_I2077 (.Y(N7767), .A(N7381), .B(N7467));
AO21XL inst_cellmath__198_0_I2078 (.Y(N7917), .A0(N7668), .A1(N7612), .B0(N7528));
AND2XL inst_cellmath__198_0_I2079 (.Y(N7403), .A(N7668), .B(N7747));
AO21XL inst_cellmath__198_0_I2080 (.Y(N7551), .A0(N7302), .A1(N7892), .B0(N7807));
AND2XL inst_cellmath__198_0_I2081 (.Y(N7689), .A(N7302), .B(N7381));
AO21XL inst_cellmath__198_0_I2082 (.Y(N7299), .A0(N7703), .A1(N7605), .B0(N7561));
AO21XL inst_cellmath__198_0_I2083 (.Y(N7584), .A0(N7338), .A1(N7627), .B0(N7842));
AO21XL inst_cellmath__198_0_I2084 (.Y(N7863), .A0(N7624), .A1(N7644), .B0(N7481));
AO21XL inst_cellmath__198_0_I2085 (.Y(N7502), .A0(N7907), .A1(N7932), .B0(N7758));
AO21XL inst_cellmath__198_0_I2086 (.Y(N7779), .A0(N7541), .A1(N7561), .B0(N7393));
AND2XL inst_cellmath__198_0_I2087 (.Y(N7929), .A(N7541), .B(N7703));
AO21XL inst_cellmath__198_0_I2088 (.Y(N7416), .A0(N7820), .A1(N7842), .B0(N7681));
AND2XL inst_cellmath__198_0_I2089 (.Y(N7559), .A(N7820), .B(N7338));
AO21XL inst_cellmath__198_0_I2090 (.Y(N7701), .A0(N7458), .A1(N7481), .B0(N7313));
AND2XL inst_cellmath__198_0_I2091 (.Y(N7840), .A(N7458), .B(N7624));
AO21XL inst_cellmath__198_0_I2092 (.Y(N7335), .A0(N7737), .A1(N7758), .B0(N7598));
AND2XL inst_cellmath__198_0_I2093 (.Y(N7478), .A(N7737), .B(N7907));
AO21XL inst_cellmath__198_0_I2094 (.Y(N7622), .A0(N7371), .A1(N7393), .B0(N7879));
AND2XL inst_cellmath__198_0_I2095 (.Y(N7756), .A(N7371), .B(N7541));
AO21XL inst_cellmath__198_0_I2096 (.Y(N7902), .A0(N7656), .A1(N7681), .B0(N7515));
AO21XL inst_cellmath__198_0_I2097 (.Y(N7537), .A0(N7287), .A1(N7313), .B0(N7793));
AO21XL inst_cellmath__198_0_I2098 (.Y(N7816), .A0(N7573), .A1(N7598), .B0(N7429));
AO21XL inst_cellmath__198_0_I2099 (.Y(N7454), .A0(N7850), .A1(N7879), .B0(N7714));
AND2XL inst_cellmath__198_0_I2100 (.Y(N7594), .A(N7850), .B(N7371));
AO21XL inst_cellmath__198_0_I2101 (.Y(N7733), .A0(N7489), .A1(N7515), .B0(N7348));
AND2XL inst_cellmath__198_0_I2102 (.Y(N7874), .A(N7489), .B(N7656));
AO21XL inst_cellmath__198_0_I2103 (.Y(N7368), .A0(N7767), .A1(N7793), .B0(N7634));
AND2XL inst_cellmath__198_0_I2104 (.Y(N7511), .A(N7767), .B(N7287));
AO21XL inst_cellmath__198_0_I2105 (.Y(N7652), .A0(N7403), .A1(N7429), .B0(N7917));
AND2XL inst_cellmath__198_0_I2106 (.Y(N7789), .A(N7403), .B(N7573));
AO21XL inst_cellmath__198_0_I2107 (.Y(N7939), .A0(N7689), .A1(N7714), .B0(N7551));
AND2XL inst_cellmath__198_0_I2108 (.Y(N7425), .A(N7689), .B(N7850));
AO21XL inst_cellmath__198_0_I2109 (.Y(N7836), .A0(N7594), .A1(N7779), .B0(N7454));
AND2XL inst_cellmath__198_0_I2110 (.Y(N7331), .A(N7594), .B(N7929));
AO21XL inst_cellmath__198_0_I2111 (.Y(N7472), .A0(N7874), .A1(N7416), .B0(N7733));
AND2XL inst_cellmath__198_0_I2112 (.Y(N7617), .A(N7874), .B(N7559));
AO21XL inst_cellmath__198_0_I2113 (.Y(N7752), .A0(N7511), .A1(N7701), .B0(N7368));
AND2XL inst_cellmath__198_0_I2114 (.Y(N7897), .A(N7511), .B(N7840));
AO21XL inst_cellmath__198_0_I2115 (.Y(N7387), .A0(N7789), .A1(N7335), .B0(N7652));
AND2XL inst_cellmath__198_0_I2116 (.Y(N7533), .A(N7789), .B(N7478));
AO21XL inst_cellmath__198_0_I2117 (.Y(N7674), .A0(N7425), .A1(N7622), .B0(N7939));
AND2XL inst_cellmath__198_0_I2118 (.Y(N7812), .A(N7425), .B(N7756));
AOI21XL inst_cellmath__198_0_I2119 (.Y(N7798), .A0(N7929), .A1(N7605), .B0(N7779));
AOI21XL inst_cellmath__198_0_I2120 (.Y(N7295), .A0(N7559), .A1(N7627), .B0(N7416));
AOI21XL inst_cellmath__198_0_I2121 (.Y(N7435), .A0(N7840), .A1(N7644), .B0(N7701));
AOI21XL inst_cellmath__198_0_I2122 (.Y(N7579), .A0(N7478), .A1(N7932), .B0(N7335));
AOI21XL inst_cellmath__198_0_I2123 (.Y(N7721), .A0(N7756), .A1(N7299), .B0(N7622));
AOI31X1 inst_cellmath__198_0_I2124 (.Y(N7857), .A0(N7656), .A1(N7820), .A2(N7584), .B0(N7902));
AOI31X1 inst_cellmath__198_0_I2125 (.Y(N7352), .A0(N7287), .A1(N7458), .A2(N7863), .B0(N7537));
AOI31X1 inst_cellmath__198_0_I2126 (.Y(N7498), .A0(N7573), .A1(N7737), .A2(N7502), .B0(N7816));
AO21XL inst_cellmath__198_0_I2127 (.Y(N7578), .A0(N7331), .A1(N7605), .B0(N7836));
AO21XL inst_cellmath__198_0_I2128 (.Y(N7855), .A0(N7617), .A1(N7627), .B0(N7472));
AO21XL inst_cellmath__198_0_I2129 (.Y(N7496), .A0(N7897), .A1(N7644), .B0(N7752));
AO21XL inst_cellmath__198_0_I2130 (.Y(N7773), .A0(N7533), .A1(N7932), .B0(N7387));
AO21XL inst_cellmath__198_0_I2131 (.Y(N7409), .A0(N7812), .A1(N7299), .B0(N7674));
NAND2BXL inst_cellmath__198_0_I2137 (.Y(N7564), .AN(N7353), .B(N7497));
NAND2BXL inst_cellmath__198_0_I2138 (.Y(N7340), .AN(N7638), .B(N7774));
NAND2BXL inst_cellmath__198_0_I2139 (.Y(N7760), .AN(N7923), .B(N7410));
NAND2BXL inst_cellmath__198_0_I2140 (.Y(N7542), .AN(N7555), .B(N7696));
NAND2BXL inst_cellmath__198_0_I2141 (.Y(N7315), .AN(N7833), .B(N7329));
NAND2BXL inst_cellmath__198_0_I2142 (.Y(N7738), .AN(N7470), .B(N7615));
NAND2BXL inst_cellmath__198_0_I2143 (.Y(N7516), .AN(N7750), .B(N7895));
NAND2BXL inst_cellmath__198_0_I2144 (.Y(N7289), .AN(N7385), .B(N7531));
NAND2BXL inst_cellmath__198_0_I2145 (.Y(N7715), .AN(N7671), .B(N7810));
NAND2BXL inst_cellmath__198_0_I2146 (.Y(N7491), .AN(N7305), .B(N7447));
NAND2BXL inst_cellmath__198_0_I2147 (.Y(N7919), .AN(N7590), .B(N7728));
NAND2BXL inst_cellmath__198_0_I2148 (.Y(N7691), .AN(N7868), .B(N7362));
NAND2BXL inst_cellmath__198_0_I2149 (.Y(N7466), .AN(N7506), .B(N7646));
NAND2BXL inst_cellmath__198_0_I2150 (.Y(N7890), .AN(N7784), .B(N7934));
NAND2BXL inst_cellmath__198_0_I2151 (.Y(N7666), .AN(N7420), .B(N7566));
NOR2BX1 inst_cellmath__198_0_I2152 (.Y(N7443), .AN(N7940), .B(N7427));
XOR2XL inst_cellmath__198_0_I2159 (.Y(inst_cellmath__198[18]), .A(N7863), .B(N7340));
XOR2XL inst_cellmath__198_0_I2160 (.Y(inst_cellmath__198[19]), .A(N7502), .B(N7760));
XNOR2X1 inst_cellmath__198_0_I2161 (.Y(inst_cellmath__198[20]), .A(N7798), .B(N7542));
XNOR2X1 inst_cellmath__198_0_I2162 (.Y(inst_cellmath__198[21]), .A(N7295), .B(N7315));
XNOR2X1 inst_cellmath__198_0_I2163 (.Y(inst_cellmath__198[22]), .A(N7435), .B(N7738));
XNOR2X1 inst_cellmath__198_0_I2164 (.Y(inst_cellmath__198[23]), .A(N7579), .B(N7516));
XNOR2X1 inst_cellmath__198_0_I2165 (.Y(inst_cellmath__198[24]), .A(N7721), .B(N7289));
XNOR2X1 inst_cellmath__198_0_I2166 (.Y(inst_cellmath__198[25]), .A(N7857), .B(N7715));
XNOR2X1 inst_cellmath__198_0_I2167 (.Y(inst_cellmath__198[26]), .A(N7352), .B(N7491));
XNOR2X1 inst_cellmath__198_0_I2168 (.Y(inst_cellmath__198[27]), .A(N7498), .B(N7919));
XOR2XL inst_cellmath__198_0_I2169 (.Y(inst_cellmath__198[28]), .A(N7578), .B(N7691));
XOR2XL inst_cellmath__198_0_I2170 (.Y(inst_cellmath__198[29]), .A(N7855), .B(N7466));
XOR2XL inst_cellmath__198_0_I2171 (.Y(inst_cellmath__198[30]), .A(N7496), .B(N7890));
XOR2XL inst_cellmath__198_0_I2172 (.Y(inst_cellmath__198[31]), .A(N7773), .B(N7666));
XOR2XL inst_cellmath__198_0_I2173 (.Y(inst_cellmath__198[32]), .A(N7409), .B(N7443));
INVXL inst_cellmath__203_0_I2174 (.Y(N10240), .A(inst_cellmath__197[0]));
INVXL inst_cellmath__203_0_I2175 (.Y(N8905), .A(inst_cellmath__197[1]));
INVXL inst_cellmath__203_0_I2176 (.Y(N9281), .A(inst_cellmath__197[2]));
INVXL inst_cellmath__203_0_I2177 (.Y(N9673), .A(inst_cellmath__197[3]));
INVXL inst_cellmath__203_0_I2178 (.Y(N10037), .A(inst_cellmath__197[4]));
INVXL inst_cellmath__203_0_I2179 (.Y(N8704), .A(inst_cellmath__197[5]));
INVXL inst_cellmath__203_0_I2180 (.Y(N9054), .A(inst_cellmath__197[6]));
INVXL inst_cellmath__203_0_I2181 (.Y(N9446), .A(inst_cellmath__197[7]));
INVXL inst_cellmath__203_0_I2182 (.Y(N9822), .A(inst_cellmath__197[8]));
INVXL inst_cellmath__203_0_I2183 (.Y(N10184), .A(inst_cellmath__197[9]));
INVXL inst_cellmath__203_0_I2184 (.Y(N8844), .A(inst_cellmath__197[10]));
INVXL inst_cellmath__203_0_I2185 (.Y(N9213), .A(inst_cellmath__197[11]));
INVXL inst_cellmath__203_0_I2186 (.Y(N9605), .A(inst_cellmath__197[12]));
INVXL inst_cellmath__203_0_I2187 (.Y(N9973), .A(inst_cellmath__197[13]));
INVXL inst_cellmath__203_0_I2188 (.Y(N8654), .A(inst_cellmath__197[14]));
INVXL inst_cellmath__203_0_I2189 (.Y(N8994), .A(inst_cellmath__197[15]));
INVXL inst_cellmath__203_0_I2190 (.Y(N9376), .A(inst_cellmath__197[16]));
INVXL inst_cellmath__203_0_I2191 (.Y(N9760), .A(inst_cellmath__197[17]));
INVXL inst_cellmath__203_0_I2192 (.Y(N10120), .A(inst_cellmath__197[18]));
INVXL inst_cellmath__203_0_I2193 (.Y(N8781), .A(inst_cellmath__197[19]));
XNOR2X1 inst_cellmath__203_0_I8338 (.Y(N9147), .A(N7584), .B(N7564));
NOR2XL inst_cellmath__203_0_I2196 (.Y(N10207), .A(N9147), .B(N8905));
NOR2XL inst_cellmath__203_0_I2197 (.Y(N9240), .A(N9147), .B(N9281));
NOR2XL inst_cellmath__203_0_I2198 (.Y(N9998), .A(N9147), .B(N9673));
NOR2XL inst_cellmath__203_0_I2199 (.Y(N9014), .A(N9147), .B(N10037));
NOR2XL inst_cellmath__203_0_I2200 (.Y(N9787), .A(N9147), .B(N8704));
NOR2XL inst_cellmath__203_0_I2201 (.Y(N8804), .A(N9147), .B(N9054));
NOR2XL inst_cellmath__203_0_I2202 (.Y(N9563), .A(N9147), .B(N9446));
NOR2XL inst_cellmath__203_0_I2203 (.Y(N8621), .A(N9147), .B(N9822));
NOR2XL inst_cellmath__203_0_I2204 (.Y(N9334), .A(N9147), .B(N10184));
NOR2XL inst_cellmath__203_0_I2205 (.Y(N10081), .A(N9147), .B(N8844));
NOR2XL inst_cellmath__203_0_I2206 (.Y(N9105), .A(N9147), .B(N9213));
NOR2XL inst_cellmath__203_0_I2207 (.Y(N9878), .A(N9147), .B(N9605));
NOR2XL inst_cellmath__203_0_I2208 (.Y(N8890), .A(N9147), .B(N9973));
NOR2XL inst_cellmath__203_0_I2209 (.Y(N9662), .A(N9147), .B(N8654));
NOR2XL inst_cellmath__203_0_I2210 (.Y(N8693), .A(N9147), .B(N8994));
NOR2XL inst_cellmath__203_0_I2211 (.Y(N9430), .A(N9147), .B(N9376));
NOR2XL inst_cellmath__203_0_I2212 (.Y(N10174), .A(N9147), .B(N9760));
NOR2XL inst_cellmath__203_0_I2213 (.Y(N9201), .A(N9147), .B(N10120));
NOR2XL inst_cellmath__203_0_I2214 (.Y(N9963), .A(N9147), .B(N8781));
INVXL inst_cellmath__203_0_I2215 (.Y(N8599), .A(inst_cellmath__198[18]));
NAND2BX1 inst_cellmath__203_0_I2216 (.Y(N8931), .AN(inst_cellmath__198[19]), .B(inst_cellmath__198[18]));
INVXL inst_cellmath__203_0_I2217 (.Y(N9310), .A(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I2218 (.Y(N9632), .A(N10240), .B(N8599));
MXI2XL inst_cellmath__203_0_I2219 (.Y(inst_cellmath__203__W0[1]), .A(N9310), .B(N8931), .S0(N9632));
MXI2XL inst_cellmath__203_0_I2220 (.Y(N9565), .A(N8905), .B(N10240), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2221 (.Y(N9295), .A(N9310), .B(N8931), .S0(N9565));
MXI2XL inst_cellmath__203_0_I2222 (.Y(N9498), .A(N9281), .B(N8905), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2223 (.Y(N9687), .A(N9310), .B(N8931), .S0(N9498));
MXI2XL inst_cellmath__203_0_I2224 (.Y(N9433), .A(N9673), .B(N9281), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2225 (.Y(N10051), .A(N9310), .B(N8931), .S0(N9433));
MXI2XL inst_cellmath__203_0_I2226 (.Y(N9365), .A(N10037), .B(N9673), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2227 (.Y(N8716), .A(N9310), .B(N8931), .S0(N9365));
MXI2XL inst_cellmath__203_0_I2228 (.Y(N9298), .A(N8704), .B(N10037), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2229 (.Y(N9068), .A(N9310), .B(N8931), .S0(N9298));
MXI2XL inst_cellmath__203_0_I2230 (.Y(N9233), .A(N9054), .B(N8704), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2231 (.Y(N9461), .A(N9310), .B(N8931), .S0(N9233));
MXI2XL inst_cellmath__203_0_I2232 (.Y(N9168), .A(N9446), .B(N9054), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2233 (.Y(N9840), .A(N9310), .B(N8931), .S0(N9168));
MXI2XL inst_cellmath__203_0_I2234 (.Y(N9099), .A(N9822), .B(N9446), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2235 (.Y(N10198), .A(N9310), .B(N8931), .S0(N9099));
MXI2XL inst_cellmath__203_0_I2236 (.Y(N9033), .A(N10184), .B(N9822), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2237 (.Y(N8858), .A(N9310), .B(N8931), .S0(N9033));
MXI2XL inst_cellmath__203_0_I2238 (.Y(N8976), .A(N8844), .B(N10184), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2239 (.Y(N9229), .A(N9310), .B(N8931), .S0(N8976));
MXI2XL inst_cellmath__203_0_I2240 (.Y(N8913), .A(N9213), .B(N8844), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2241 (.Y(N9622), .A(N9310), .B(N8931), .S0(N8913));
MXI2XL inst_cellmath__203_0_I2242 (.Y(N8853), .A(N9605), .B(N9213), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2243 (.Y(N9989), .A(N9310), .B(N8931), .S0(N8853));
MXI2XL inst_cellmath__203_0_I2244 (.Y(N8792), .A(N9973), .B(N9605), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2245 (.Y(N8666), .A(N9310), .B(N8931), .S0(N8792));
MXI2XL inst_cellmath__203_0_I2246 (.Y(N8735), .A(N8654), .B(N9973), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2247 (.Y(N9006), .A(N9310), .B(N8931), .S0(N8735));
MXI2XL inst_cellmath__203_0_I2248 (.Y(N8681), .A(N8994), .B(N8654), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2249 (.Y(N9393), .A(N9310), .B(N8931), .S0(N8681));
MXI2XL inst_cellmath__203_0_I2250 (.Y(N8634), .A(N9376), .B(N8994), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2251 (.Y(N9779), .A(N9310), .B(N8931), .S0(N8634));
MXI2XL inst_cellmath__203_0_I2252 (.Y(N8582), .A(N9760), .B(N9376), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2253 (.Y(N10136), .A(N9310), .B(N8931), .S0(N8582));
MXI2XL inst_cellmath__203_0_I2254 (.Y(N10188), .A(N10120), .B(N9760), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2255 (.Y(N8798), .A(N9310), .B(N8931), .S0(N10188));
MXI2XL inst_cellmath__203_0_I2256 (.Y(N10125), .A(N8781), .B(N10120), .S0(N8599));
MXI2XL inst_cellmath__203_0_I2257 (.Y(N9164), .A(N9310), .B(N8931), .S0(N10125));
NAND2XL inst_cellmath__203_0_I2258 (.Y(N10062), .A(N8781), .B(N8599));
MXI2XL inst_cellmath__203_0_I2259 (.Y(N9556), .A(N9310), .B(N8931), .S0(N10062));
XNOR2X1 inst_cellmath__203_0_I2260 (.Y(N9331), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I2261 (.Y(N9021), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
OAI2BB1X1 inst_cellmath__203_0_I2262 (.Y(N8947), .A0N(inst_cellmath__198[20]), .A1N(inst_cellmath__198[19]), .B0(inst_cellmath__198[21]));
INVXL inst_cellmath__203_0_I2263 (.Y(N9696), .A(N8947));
OR2XL inst_cellmath__203_0_I2264 (.Y(N9082), .A(N9021), .B(inst_cellmath__198[21]));
INVXL inst_cellmath__203_0_I2265 (.Y(N9474), .A(N9696));
NOR2XL inst_cellmath__203_0_I2266 (.Y(N9729), .A(N10240), .B(N9331));
MXI2XL inst_cellmath__203_0_I2267 (.Y(N9871), .A(N9474), .B(N9082), .S0(N9729));
MXI2XL inst_cellmath__203_0_I2268 (.Y(N9669), .A(N8905), .B(N10240), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2269 (.Y(N10222), .A(N9474), .B(N9082), .S0(N9669));
MXI2XL inst_cellmath__203_0_I2270 (.Y(N9601), .A(N9281), .B(N8905), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2271 (.Y(N8882), .A(N9474), .B(N9082), .S0(N9601));
MXI2XL inst_cellmath__203_0_I2272 (.Y(N9534), .A(N9673), .B(N9281), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2273 (.Y(N9263), .A(N9474), .B(N9082), .S0(N9534));
MXI2XL inst_cellmath__203_0_I2274 (.Y(N9471), .A(N10037), .B(N9673), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2275 (.Y(N9653), .A(N9474), .B(N9082), .S0(N9471));
MXI2XL inst_cellmath__203_0_I2276 (.Y(N9400), .A(N8704), .B(N10037), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2277 (.Y(N10017), .A(N9474), .B(N9082), .S0(N9400));
MXI2XL inst_cellmath__203_0_I2278 (.Y(N9335), .A(N9054), .B(N8704), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2279 (.Y(N8687), .A(N9474), .B(N9082), .S0(N9335));
MXI2XL inst_cellmath__203_0_I2280 (.Y(N9268), .A(N9446), .B(N9054), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2281 (.Y(N9032), .A(N9474), .B(N9082), .S0(N9268));
MXI2XL inst_cellmath__203_0_I2282 (.Y(N9202), .A(N9822), .B(N9446), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2283 (.Y(N9423), .A(N9474), .B(N9082), .S0(N9202));
MXI2XL inst_cellmath__203_0_I2284 (.Y(N9132), .A(N10184), .B(N9822), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2285 (.Y(N9807), .A(N9474), .B(N9082), .S0(N9132));
MXI2XL inst_cellmath__203_0_I2286 (.Y(N9069), .A(N8844), .B(N10184), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2287 (.Y(N10165), .A(N9474), .B(N9082), .S0(N9069));
MXI2XL inst_cellmath__203_0_I2288 (.Y(N9007), .A(N9213), .B(N8844), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2289 (.Y(N8823), .A(N9474), .B(N9082), .S0(N9007));
MXI2XL inst_cellmath__203_0_I2290 (.Y(N8948), .A(N9605), .B(N9213), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2291 (.Y(N9196), .A(N9474), .B(N9082), .S0(N8948));
MXI2XL inst_cellmath__203_0_I2292 (.Y(N8883), .A(N9973), .B(N9605), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2293 (.Y(N9589), .A(N9474), .B(N9082), .S0(N8883));
MXI2XL inst_cellmath__203_0_I2294 (.Y(N8824), .A(N8654), .B(N9973), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2295 (.Y(N9954), .A(N9474), .B(N9082), .S0(N8824));
MXI2XL inst_cellmath__203_0_I2296 (.Y(N8764), .A(N8994), .B(N8654), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2297 (.Y(N8639), .A(N9474), .B(N9082), .S0(N8764));
MXI2XL inst_cellmath__203_0_I2298 (.Y(N8711), .A(N9376), .B(N8994), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2299 (.Y(N8975), .A(N9474), .B(N9082), .S0(N8711));
MXI2XL inst_cellmath__203_0_I2300 (.Y(N8660), .A(N9760), .B(N9376), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2301 (.Y(N9356), .A(N9474), .B(N9082), .S0(N8660));
MXI2XL inst_cellmath__203_0_I2302 (.Y(N8607), .A(N10120), .B(N9760), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2303 (.Y(N9743), .A(N9474), .B(N9082), .S0(N8607));
MXI2XL inst_cellmath__203_0_I2304 (.Y(N10215), .A(N8781), .B(N10120), .S0(N9331));
MXI2XL inst_cellmath__203_0_I2305 (.Y(N10101), .A(N9474), .B(N9082), .S0(N10215));
NAND2XL inst_cellmath__203_0_I2306 (.Y(N10157), .A(N8781), .B(N9331));
MXI2XL inst_cellmath__203_0_I2307 (.Y(N8763), .A(N9474), .B(N9082), .S0(N10157));
XNOR2X1 inst_cellmath__203_0_I2308 (.Y(N8586), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
NOR2XL inst_cellmath__203_0_I2309 (.Y(N9121), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
OAI2BB1X1 inst_cellmath__203_0_I2310 (.Y(N9895), .A0N(inst_cellmath__198[22]), .A1N(inst_cellmath__198[21]), .B0(inst_cellmath__198[23]));
INVXL inst_cellmath__203_0_I2311 (.Y(N9853), .A(N9895));
OR2XL inst_cellmath__203_0_I2312 (.Y(N9246), .A(N9121), .B(inst_cellmath__198[23]));
INVXL inst_cellmath__203_0_I2313 (.Y(N9634), .A(N9853));
NOR2XL inst_cellmath__203_0_I2314 (.Y(N9823), .A(N10240), .B(N8586));
MXI2XL inst_cellmath__203_0_I2315 (.Y(N9062), .A(N9634), .B(N9246), .S0(N9823));
MXI2XL inst_cellmath__203_0_I2316 (.Y(N9762), .A(N8905), .B(N10240), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2317 (.Y(N9456), .A(N9634), .B(N9246), .S0(N9762));
MXI2XL inst_cellmath__203_0_I2318 (.Y(N9698), .A(N9281), .B(N8905), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2319 (.Y(N9831), .A(N9634), .B(N9246), .S0(N9698));
MXI2XL inst_cellmath__203_0_I2320 (.Y(N9636), .A(N9673), .B(N9281), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2321 (.Y(N10191), .A(N9634), .B(N9246), .S0(N9636));
MXI2XL inst_cellmath__203_0_I2322 (.Y(N9569), .A(N10037), .B(N9673), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2323 (.Y(N8851), .A(N9634), .B(N9246), .S0(N9569));
MXI2XL inst_cellmath__203_0_I2324 (.Y(N9501), .A(N8704), .B(N10037), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2325 (.Y(N9222), .A(N9634), .B(N9246), .S0(N9501));
MXI2XL inst_cellmath__203_0_I2326 (.Y(N9437), .A(N9054), .B(N8704), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2327 (.Y(N9614), .A(N9634), .B(N9246), .S0(N9437));
MXI2XL inst_cellmath__203_0_I2328 (.Y(N9368), .A(N9446), .B(N9054), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2329 (.Y(N9981), .A(N9634), .B(N9246), .S0(N9368));
MXI2XL inst_cellmath__203_0_I2330 (.Y(N9301), .A(N9822), .B(N9446), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2331 (.Y(N8659), .A(N9634), .B(N9246), .S0(N9301));
MXI2XL inst_cellmath__203_0_I2332 (.Y(N9239), .A(N10184), .B(N9822), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2333 (.Y(N9001), .A(N9634), .B(N9246), .S0(N9239));
MXI2XL inst_cellmath__203_0_I2334 (.Y(N9172), .A(N8844), .B(N10184), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2335 (.Y(N9387), .A(N9634), .B(N9246), .S0(N9172));
MXI2XL inst_cellmath__203_0_I2336 (.Y(N9102), .A(N9213), .B(N8844), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2337 (.Y(N9770), .A(N9634), .B(N9246), .S0(N9102));
MXI2XL inst_cellmath__203_0_I2338 (.Y(N9038), .A(N9605), .B(N9213), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2339 (.Y(N10129), .A(N9634), .B(N9246), .S0(N9038));
MXI2XL inst_cellmath__203_0_I2340 (.Y(N8980), .A(N9973), .B(N9605), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2341 (.Y(N8790), .A(N9634), .B(N9246), .S0(N8980));
MXI2XL inst_cellmath__203_0_I2342 (.Y(N8917), .A(N8654), .B(N9973), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2343 (.Y(N9156), .A(N9634), .B(N9246), .S0(N8917));
MXI2XL inst_cellmath__203_0_I2344 (.Y(N8856), .A(N8994), .B(N8654), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2345 (.Y(N9547), .A(N9634), .B(N9246), .S0(N8856));
MXI2XL inst_cellmath__203_0_I2346 (.Y(N8795), .A(N9376), .B(N8994), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2347 (.Y(N9921), .A(N9634), .B(N9246), .S0(N8795));
MXI2XL inst_cellmath__203_0_I2348 (.Y(N8739), .A(N9760), .B(N9376), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2349 (.Y(N8606), .A(N9634), .B(N9246), .S0(N8739));
MXI2XL inst_cellmath__203_0_I2350 (.Y(N8685), .A(N10120), .B(N9760), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2351 (.Y(N8941), .A(N9634), .B(N9246), .S0(N8685));
MXI2XL inst_cellmath__203_0_I2352 (.Y(N8637), .A(N8781), .B(N10120), .S0(N8586));
MXI2XL inst_cellmath__203_0_I2353 (.Y(N9322), .A(N9634), .B(N9246), .S0(N8637));
NAND2XL inst_cellmath__203_0_I2354 (.Y(N8585), .A(N8781), .B(N8586));
MXI2XL inst_cellmath__203_0_I2355 (.Y(N9706), .A(N9634), .B(N9246), .S0(N8585));
XNOR2X1 inst_cellmath__203_0_I2356 (.Y(N9483), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
NOR2XL inst_cellmath__203_0_I2357 (.Y(N9220), .A(inst_cellmath__198[24]), .B(inst_cellmath__198[23]));
OAI2BB1X1 inst_cellmath__203_0_I2358 (.Y(N9090), .A0N(inst_cellmath__198[24]), .A1N(inst_cellmath__198[23]), .B0(inst_cellmath__198[25]));
INVXL inst_cellmath__203_0_I2359 (.Y(N10000), .A(N9090));
OR2XL inst_cellmath__203_0_I2360 (.Y(N9404), .A(N9220), .B(inst_cellmath__198[25]));
INVXL inst_cellmath__203_0_I2361 (.Y(N9789), .A(N10000));
NOR2XL inst_cellmath__203_0_I2362 (.Y(N9918), .A(N10240), .B(N9483));
MXI2XL inst_cellmath__203_0_I2363 (.Y(N10007), .A(N9789), .B(N9404), .S0(N9918));
MXI2XL inst_cellmath__203_0_I2364 (.Y(N9860), .A(N8905), .B(N10240), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2365 (.Y(N8679), .A(N9789), .B(N9404), .S0(N9860));
MXI2XL inst_cellmath__203_0_I2366 (.Y(N9796), .A(N9281), .B(N8905), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2367 (.Y(N9026), .A(N9789), .B(N9404), .S0(N9796));
MXI2XL inst_cellmath__203_0_I2368 (.Y(N9732), .A(N9673), .B(N9281), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2369 (.Y(N9414), .A(N9789), .B(N9404), .S0(N9732));
MXI2XL inst_cellmath__203_0_I2370 (.Y(N9672), .A(N10037), .B(N9673), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2371 (.Y(N9798), .A(N9789), .B(N9404), .S0(N9672));
MXI2XL inst_cellmath__203_0_I2372 (.Y(N9604), .A(N8704), .B(N10037), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2373 (.Y(N10156), .A(N9789), .B(N9404), .S0(N9604));
MXI2XL inst_cellmath__203_0_I2374 (.Y(N9536), .A(N9054), .B(N8704), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2375 (.Y(N8816), .A(N9789), .B(N9404), .S0(N9536));
MXI2XL inst_cellmath__203_0_I2376 (.Y(N9473), .A(N9446), .B(N9054), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2377 (.Y(N9187), .A(N9789), .B(N9404), .S0(N9473));
MXI2XL inst_cellmath__203_0_I2378 (.Y(N9403), .A(N9822), .B(N9446), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2379 (.Y(N9577), .A(N9789), .B(N9404), .S0(N9403));
MXI2XL inst_cellmath__203_0_I2380 (.Y(N9338), .A(N10184), .B(N9822), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2381 (.Y(N9945), .A(N9789), .B(N9404), .S0(N9338));
MXI2XL inst_cellmath__203_0_I2382 (.Y(N9271), .A(N8844), .B(N10184), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2383 (.Y(N8630), .A(N9789), .B(N9404), .S0(N9271));
MXI2XL inst_cellmath__203_0_I2384 (.Y(N9204), .A(N9213), .B(N8844), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2385 (.Y(N8966), .A(N9789), .B(N9404), .S0(N9204));
MXI2XL inst_cellmath__203_0_I2386 (.Y(N9134), .A(N9605), .B(N9213), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2387 (.Y(N9348), .A(N9789), .B(N9404), .S0(N9134));
MXI2XL inst_cellmath__203_0_I2388 (.Y(N9071), .A(N9973), .B(N9605), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2389 (.Y(N9733), .A(N9789), .B(N9404), .S0(N9071));
MXI2XL inst_cellmath__203_0_I2390 (.Y(N9010), .A(N8654), .B(N9973), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2391 (.Y(N10093), .A(N9789), .B(N9404), .S0(N9010));
MXI2XL inst_cellmath__203_0_I2392 (.Y(N8951), .A(N8994), .B(N8654), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2393 (.Y(N8757), .A(N9789), .B(N9404), .S0(N8951));
MXI2XL inst_cellmath__203_0_I2394 (.Y(N8884), .A(N9376), .B(N8994), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2395 (.Y(N9120), .A(N9789), .B(N9404), .S0(N8884));
MXI2XL inst_cellmath__203_0_I2396 (.Y(N8828), .A(N9760), .B(N9376), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2397 (.Y(N9509), .A(N9789), .B(N9404), .S0(N8828));
MXI2XL inst_cellmath__203_0_I2398 (.Y(N8767), .A(N10120), .B(N9760), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2399 (.Y(N9888), .A(N9789), .B(N9404), .S0(N8767));
MXI2XL inst_cellmath__203_0_I2400 (.Y(N8712), .A(N8781), .B(N10120), .S0(N9483));
MXI2XL inst_cellmath__203_0_I2401 (.Y(N8580), .A(N9789), .B(N9404), .S0(N8712));
NAND2XL inst_cellmath__203_0_I2402 (.Y(N8664), .A(N8781), .B(N9483));
MXI2XL inst_cellmath__203_0_I2403 (.Y(N8906), .A(N9789), .B(N9404), .S0(N8664));
XNOR2X1 inst_cellmath__203_0_I2404 (.Y(N8705), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NOR2XL inst_cellmath__203_0_I2405 (.Y(N9325), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
OAI2BB1X1 inst_cellmath__203_0_I2406 (.Y(N10039), .A0N(inst_cellmath__198[26]), .A1N(inst_cellmath__198[25]), .B0(inst_cellmath__198[27]));
INVXL inst_cellmath__203_0_I2407 (.Y(N10148), .A(N10039));
OR2XL inst_cellmath__203_0_I2408 (.Y(N9567), .A(N9325), .B(inst_cellmath__198[27]));
INVXL inst_cellmath__203_0_I2409 (.Y(N9938), .A(N10148));
NOR2XL inst_cellmath__203_0_I2410 (.Y(N10010), .A(N10240), .B(N8705));
MXI2XL inst_cellmath__203_0_I2411 (.Y(N9214), .A(N9938), .B(N9567), .S0(N10010));
MXI2XL inst_cellmath__203_0_I2412 (.Y(N9949), .A(N8905), .B(N10240), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2413 (.Y(N9606), .A(N9938), .B(N9567), .S0(N9949));
MXI2XL inst_cellmath__203_0_I2414 (.Y(N9890), .A(N9281), .B(N8905), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2415 (.Y(N9975), .A(N9938), .B(N9567), .S0(N9890));
MXI2XL inst_cellmath__203_0_I2416 (.Y(N9826), .A(N9673), .B(N9281), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2417 (.Y(N8655), .A(N9938), .B(N9567), .S0(N9826));
MXI2XL inst_cellmath__203_0_I2418 (.Y(N9765), .A(N10037), .B(N9673), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2419 (.Y(N8996), .A(N9938), .B(N9567), .S0(N9765));
MXI2XL inst_cellmath__203_0_I2420 (.Y(N9700), .A(N8704), .B(N10037), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2421 (.Y(N9377), .A(N9938), .B(N9567), .S0(N9700));
MXI2XL inst_cellmath__203_0_I2422 (.Y(N9640), .A(N9054), .B(N8704), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2423 (.Y(N9761), .A(N9938), .B(N9567), .S0(N9640));
MXI2XL inst_cellmath__203_0_I2424 (.Y(N9573), .A(N9446), .B(N9054), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2425 (.Y(N10122), .A(N9938), .B(N9567), .S0(N9573));
MXI2XL inst_cellmath__203_0_I2426 (.Y(N9505), .A(N9822), .B(N9446), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2427 (.Y(N8783), .A(N9938), .B(N9567), .S0(N9505));
MXI2XL inst_cellmath__203_0_I2428 (.Y(N9442), .A(N10184), .B(N9822), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2429 (.Y(N9148), .A(N9938), .B(N9567), .S0(N9442));
MXI2XL inst_cellmath__203_0_I2430 (.Y(N9372), .A(N8844), .B(N10184), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2431 (.Y(N9537), .A(N9938), .B(N9567), .S0(N9372));
MXI2XL inst_cellmath__203_0_I2432 (.Y(N9307), .A(N9213), .B(N8844), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2433 (.Y(N9913), .A(N9938), .B(N9567), .S0(N9307));
MXI2XL inst_cellmath__203_0_I2434 (.Y(N9243), .A(N9605), .B(N9213), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2435 (.Y(N8600), .A(N9938), .B(N9567), .S0(N9243));
MXI2XL inst_cellmath__203_0_I2436 (.Y(N9174), .A(N9973), .B(N9605), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2437 (.Y(N8933), .A(N9938), .B(N9567), .S0(N9174));
MXI2XL inst_cellmath__203_0_I2438 (.Y(N9106), .A(N8654), .B(N9973), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2439 (.Y(N9312), .A(N9938), .B(N9567), .S0(N9106));
MXI2XL inst_cellmath__203_0_I2440 (.Y(N9041), .A(N8994), .B(N8654), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2441 (.Y(N9697), .A(N9938), .B(N9567), .S0(N9041));
MXI2XL inst_cellmath__203_0_I2442 (.Y(N8983), .A(N9376), .B(N8994), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2443 (.Y(N10060), .A(N9938), .B(N9567), .S0(N8983));
MXI2XL inst_cellmath__203_0_I2444 (.Y(N8920), .A(N9760), .B(N9376), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2445 (.Y(N8727), .A(N9938), .B(N9567), .S0(N8920));
MXI2XL inst_cellmath__203_0_I2446 (.Y(N8859), .A(N10120), .B(N9760), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2447 (.Y(N9083), .A(N9938), .B(N9567), .S0(N8859));
MXI2XL inst_cellmath__203_0_I2448 (.Y(N8799), .A(N8781), .B(N10120), .S0(N8705));
MXI2XL inst_cellmath__203_0_I2449 (.Y(N9475), .A(N9938), .B(N9567), .S0(N8799));
NAND2XL inst_cellmath__203_0_I2450 (.Y(N8741), .A(N8781), .B(N8705));
MXI2XL inst_cellmath__203_0_I2451 (.Y(N9856), .A(N9938), .B(N9567), .S0(N8741));
XNOR2X1 inst_cellmath__203_0_I2452 (.Y(N9635), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
NOR2XL inst_cellmath__203_0_I2453 (.Y(N9424), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
OAI2BB1X1 inst_cellmath__203_0_I2454 (.Y(N9248), .A0N(inst_cellmath__198[28]), .A1N(inst_cellmath__198[27]), .B0(inst_cellmath__198[29]));
INVXL inst_cellmath__203_0_I2455 (.Y(N8623), .A(N9248));
OR2XL inst_cellmath__203_0_I2456 (.Y(N9723), .A(N9424), .B(inst_cellmath__198[29]));
INVXL inst_cellmath__203_0_I2457 (.Y(N10086), .A(N8623));
NOR2XL inst_cellmath__203_0_I2458 (.Y(N10102), .A(N10240), .B(N9635));
MXI2XL inst_cellmath__203_0_I2459 (.Y(N10149), .A(N10086), .B(N9723), .S0(N10102));
MXI2XL inst_cellmath__203_0_I2460 (.Y(N10044), .A(N8905), .B(N10240), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2461 (.Y(N8809), .A(N10086), .B(N9723), .S0(N10044));
MXI2XL inst_cellmath__203_0_I2462 (.Y(N9982), .A(N9281), .B(N8905), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2463 (.Y(N9178), .A(N10086), .B(N9723), .S0(N9982));
MXI2XL inst_cellmath__203_0_I2464 (.Y(N9922), .A(N9673), .B(N9281), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2465 (.Y(N9568), .A(N10086), .B(N9723), .S0(N9922));
MXI2XL inst_cellmath__203_0_I2466 (.Y(N9861), .A(N10037), .B(N9673), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2467 (.Y(N9939), .A(N10086), .B(N9723), .S0(N9861));
MXI2XL inst_cellmath__203_0_I2468 (.Y(N9799), .A(N8704), .B(N10037), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2469 (.Y(N8625), .A(N10086), .B(N9723), .S0(N9799));
MXI2XL inst_cellmath__203_0_I2470 (.Y(N9734), .A(N9054), .B(N8704), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2471 (.Y(N8959), .A(N10086), .B(N9723), .S0(N9734));
MXI2XL inst_cellmath__203_0_I2472 (.Y(N9675), .A(N9446), .B(N9054), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2473 (.Y(N9340), .A(N10086), .B(N9723), .S0(N9675));
MXI2XL inst_cellmath__203_0_I2474 (.Y(N9607), .A(N9822), .B(N9446), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2475 (.Y(N9726), .A(N10086), .B(N9723), .S0(N9607));
MXI2XL inst_cellmath__203_0_I2476 (.Y(N9538), .A(N10184), .B(N9822), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2477 (.Y(N10087), .A(N10086), .B(N9723), .S0(N9538));
MXI2XL inst_cellmath__203_0_I2478 (.Y(N9476), .A(N8844), .B(N10184), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2479 (.Y(N8750), .A(N10086), .B(N9723), .S0(N9476));
MXI2XL inst_cellmath__203_0_I2480 (.Y(N9406), .A(N9213), .B(N8844), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2481 (.Y(N9111), .A(N10086), .B(N9723), .S0(N9406));
MXI2XL inst_cellmath__203_0_I2482 (.Y(N9341), .A(N9605), .B(N9213), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2483 (.Y(N9500), .A(N10086), .B(N9723), .S0(N9341));
MXI2XL inst_cellmath__203_0_I2484 (.Y(N9275), .A(N9973), .B(N9605), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2485 (.Y(N9882), .A(N10086), .B(N9723), .S0(N9275));
MXI2XL inst_cellmath__203_0_I2486 (.Y(N9207), .A(N8654), .B(N9973), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2487 (.Y(N10235), .A(N10086), .B(N9723), .S0(N9207));
MXI2XL inst_cellmath__203_0_I2488 (.Y(N9139), .A(N8994), .B(N8654), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2489 (.Y(N8896), .A(N10086), .B(N9723), .S0(N9139));
MXI2XL inst_cellmath__203_0_I2490 (.Y(N9075), .A(N9376), .B(N8994), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2491 (.Y(N9274), .A(N10086), .B(N9723), .S0(N9075));
MXI2XL inst_cellmath__203_0_I2492 (.Y(N9012), .A(N9760), .B(N9376), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2493 (.Y(N9666), .A(N10086), .B(N9723), .S0(N9012));
MXI2XL inst_cellmath__203_0_I2494 (.Y(N8953), .A(N10120), .B(N9760), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2495 (.Y(N10031), .A(N10086), .B(N9723), .S0(N8953));
MXI2XL inst_cellmath__203_0_I2496 (.Y(N8889), .A(N8781), .B(N10120), .S0(N9635));
MXI2XL inst_cellmath__203_0_I2497 (.Y(N8698), .A(N10086), .B(N9723), .S0(N8889));
NAND2XL inst_cellmath__203_0_I2498 (.Y(N8832), .A(N8781), .B(N9635));
MXI2XL inst_cellmath__203_0_I2499 (.Y(N9047), .A(N10086), .B(N9723), .S0(N8832));
XNOR2X1 inst_cellmath__203_0_I2500 (.Y(N8838), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
NOR2XL inst_cellmath__203_0_I2501 (.Y(N9524), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
OAI2BB1X1 inst_cellmath__203_0_I2502 (.Y(N10180), .A0N(inst_cellmath__198[30]), .A1N(inst_cellmath__198[29]), .B0(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2503 (.Y(N8747), .A(N10180));
OR2XL inst_cellmath__203_0_I2504 (.Y(N9881), .A(N9524), .B(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2505 (.Y(N10232), .A(N8747));
NOR2XL inst_cellmath__203_0_I2506 (.Y(N10196), .A(N10240), .B(N8838));
MXI2XL inst_cellmath__203_0_I2507 (.Y(N9367), .A(N10232), .B(N9881), .S0(N10196));
MXI2XL inst_cellmath__203_0_I2508 (.Y(N10134), .A(N8905), .B(N10240), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2509 (.Y(N9755), .A(N10232), .B(N9881), .S0(N10134));
MXI2XL inst_cellmath__203_0_I2510 (.Y(N10071), .A(N9281), .B(N8905), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2511 (.Y(N10116), .A(N10232), .B(N9881), .S0(N10071));
MXI2XL inst_cellmath__203_0_I2512 (.Y(N10015), .A(N9673), .B(N9281), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2513 (.Y(N8773), .A(N10232), .B(N9881), .S0(N10015));
MXI2XL inst_cellmath__203_0_I2514 (.Y(N9953), .A(N10037), .B(N9673), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2515 (.Y(N9138), .A(N10232), .B(N9881), .S0(N9953));
MXI2XL inst_cellmath__203_0_I2516 (.Y(N9894), .A(N8704), .B(N10037), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2517 (.Y(N9531), .A(N10232), .B(N9881), .S0(N9894));
MXI2XL inst_cellmath__203_0_I2518 (.Y(N9830), .A(N9054), .B(N8704), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2519 (.Y(N9908), .A(N10232), .B(N9881), .S0(N9830));
MXI2XL inst_cellmath__203_0_I2520 (.Y(N9769), .A(N9446), .B(N9054), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2521 (.Y(N8596), .A(N10232), .B(N9881), .S0(N9769));
MXI2XL inst_cellmath__203_0_I2522 (.Y(N9705), .A(N9822), .B(N9446), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2523 (.Y(N8926), .A(N10232), .B(N9881), .S0(N9705));
MXI2XL inst_cellmath__203_0_I2524 (.Y(N9643), .A(N10184), .B(N9822), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2525 (.Y(N9304), .A(N10232), .B(N9881), .S0(N9643));
MXI2XL inst_cellmath__203_0_I2526 (.Y(N9576), .A(N8844), .B(N10184), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2527 (.Y(N9690), .A(N10232), .B(N9881), .S0(N9576));
MXI2XL inst_cellmath__203_0_I2528 (.Y(N9508), .A(N9213), .B(N8844), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2529 (.Y(N10057), .A(N10232), .B(N9881), .S0(N9508));
MXI2XL inst_cellmath__203_0_I2530 (.Y(N9445), .A(N9605), .B(N9213), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2531 (.Y(N8722), .A(N10232), .B(N9881), .S0(N9445));
MXI2XL inst_cellmath__203_0_I2532 (.Y(N9375), .A(N9973), .B(N9605), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2533 (.Y(N9074), .A(N10232), .B(N9881), .S0(N9375));
MXI2XL inst_cellmath__203_0_I2534 (.Y(N9309), .A(N8654), .B(N9973), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2535 (.Y(N9466), .A(N10232), .B(N9881), .S0(N9309));
MXI2XL inst_cellmath__203_0_I2536 (.Y(N9245), .A(N8994), .B(N8654), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2537 (.Y(N9849), .A(N10232), .B(N9881), .S0(N9245));
MXI2XL inst_cellmath__203_0_I2538 (.Y(N9176), .A(N9376), .B(N8994), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2539 (.Y(N10203), .A(N10232), .B(N9881), .S0(N9176));
MXI2XL inst_cellmath__203_0_I2540 (.Y(N9108), .A(N9760), .B(N9376), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2541 (.Y(N8863), .A(N10232), .B(N9881), .S0(N9108));
MXI2XL inst_cellmath__203_0_I2542 (.Y(N9043), .A(N10120), .B(N9760), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2543 (.Y(N9238), .A(N10232), .B(N9881), .S0(N9043));
MXI2XL inst_cellmath__203_0_I2544 (.Y(N8984), .A(N8781), .B(N10120), .S0(N8838));
MXI2XL inst_cellmath__203_0_I2545 (.Y(N9627), .A(N10232), .B(N9881), .S0(N8984));
NAND2XL inst_cellmath__203_0_I2546 (.Y(N8922), .A(N8781), .B(N8838));
MXI2XL inst_cellmath__203_0_I2547 (.Y(N9996), .A(N10232), .B(N9881), .S0(N8922));
ADDHX1 inst_cellmath__203_0_I2548 (.CO(N10143), .S(N9397), .A(inst_cellmath__198[32]), .B(inst_cellmath__198[31]));
INVXL inst_cellmath__203_0_I2549 (.Y(N8895), .A(N9397));
INVXL inst_cellmath__203_0_I2550 (.Y(N9272), .A(N10143));
NOR2XL inst_cellmath__203_0_I2551 (.Y(N10078), .A(N8895), .B(N10240));
OAI22XL inst_cellmath__203_0_I2552 (.Y(N9101), .A0(N10240), .A1(N9272), .B0(N8895), .B1(N8905));
OAI22XL inst_cellmath__203_0_I2553 (.Y(N9876), .A0(N8905), .A1(N9272), .B0(N8895), .B1(N9281));
OAI22XL inst_cellmath__203_0_I2554 (.Y(N8887), .A0(N9281), .A1(N9272), .B0(N8895), .B1(N9673));
OAI22XL inst_cellmath__203_0_I2555 (.Y(N9659), .A0(N9673), .A1(N9272), .B0(N8895), .B1(N10037));
OAI22XL inst_cellmath__203_0_I2556 (.Y(N8691), .A0(N10037), .A1(N9272), .B0(N8895), .B1(N8704));
OAI22XL inst_cellmath__203_0_I2557 (.Y(N9427), .A0(N8704), .A1(N9272), .B0(N8895), .B1(N9054));
OAI22XL inst_cellmath__203_0_I2558 (.Y(N10170), .A0(N9054), .A1(N9272), .B0(N8895), .B1(N9446));
OAI22XL inst_cellmath__203_0_I2559 (.Y(N9199), .A0(N9446), .A1(N9272), .B0(N8895), .B1(N9822));
OAI22XL inst_cellmath__203_0_I2560 (.Y(N9960), .A0(N9822), .A1(N9272), .B0(N8895), .B1(N10184));
OAI22XL inst_cellmath__203_0_I2561 (.Y(N8979), .A0(N10184), .A1(N9272), .B0(N8895), .B1(N8844));
OAI22XL inst_cellmath__203_0_I2562 (.Y(N9749), .A0(N8844), .A1(N9272), .B0(N8895), .B1(N9213));
OAI22XL inst_cellmath__203_0_I2563 (.Y(N8769), .A0(N9213), .A1(N9272), .B0(N8895), .B1(N9605));
OAI22XL inst_cellmath__203_0_I2564 (.Y(N9523), .A0(N9605), .A1(N9272), .B0(N8895), .B1(N9973));
OAI22XL inst_cellmath__203_0_I2565 (.Y(N8590), .A0(N9973), .A1(N9272), .B0(N8895), .B1(N8654));
OAI22XL inst_cellmath__203_0_I2566 (.Y(N9292), .A0(N8654), .A1(N9272), .B0(N8895), .B1(N8994));
OAI22XL inst_cellmath__203_0_I2567 (.Y(N10047), .A0(N8994), .A1(N9272), .B0(N8895), .B1(N9376));
OAI22XL inst_cellmath__203_0_I2568 (.Y(N9066), .A0(N9376), .A1(N9272), .B0(N8895), .B1(N9760));
OAI22XL inst_cellmath__203_0_I2569 (.Y(N9837), .A0(N9760), .A1(N9272), .B0(N8895), .B1(N10120));
OAI22XL inst_cellmath__203_0_I2570 (.Y(N8855), .A0(N10120), .A1(N9272), .B0(N8895), .B1(N8781));
OAI21XL inst_cellmath__203_0_I2571 (.Y(N9620), .A0(N9272), .A1(N8781), .B0(N8895));
AND2XL inst_cellmath__203_0_I2572 (.Y(N10121), .A(N9272), .B(N8895));
INVXL inst_cellmath__203_0_I2573 (.Y(N9664), .A(N742));
INVXL inst_cellmath__203_0_I2574 (.Y(N10030), .A(N743));
INVXL inst_cellmath__203_0_I2575 (.Y(N8696), .A(N744));
INVXL inst_cellmath__203_0_I2576 (.Y(N9044), .A(N745));
INVXL inst_cellmath__203_0_I2577 (.Y(N9436), .A(N746));
INVXL inst_cellmath__203_0_I2578 (.Y(N9816), .A(N747));
INVXL inst_cellmath__203_0_I2579 (.Y(N10177), .A(N748));
INVXL inst_cellmath__203_0_I2580 (.Y(N8837), .A(N749));
INVXL inst_cellmath__203_0_I2581 (.Y(N9206), .A(N750));
INVXL inst_cellmath__203_0_I2582 (.Y(N9598), .A(N751));
INVXL inst_cellmath__203_0_I2583 (.Y(N9967), .A(N752));
INVXL inst_cellmath__203_0_I2584 (.Y(N8646), .A(N753));
INVXL inst_cellmath__203_0_I2585 (.Y(N8985), .A(N754));
INVXL inst_cellmath__203_0_I2586 (.Y(N9366), .A(N755));
INVXL inst_cellmath__203_0_I2587 (.Y(N9753), .A(N756));
INVXL inst_cellmath__203_0_I2588 (.Y(N10112), .A(N757));
INVXL inst_cellmath__203_0_I2589 (.Y(N8772), .A(N758));
INVXL inst_cellmath__203_0_I2590 (.Y(N9136), .A(N759));
INVXL inst_cellmath__203_0_I2591 (.Y(N9527), .A(N760));
INVXL inst_cellmath__203_0_I2592 (.Y(N9907), .A(N761));
INVXL inst_cellmath__203_0_I2593 (.Y(N8595), .A(N762));
INVXL inst_cellmath__203_0_I2594 (.Y(N8923), .A(N763));
NOR2XL inst_cellmath__203_0_I2596 (.Y(N9492), .A(N7570), .B(N9664));
NOR2XL inst_cellmath__203_0_I2597 (.Y(N10226), .A(N7570), .B(N10030));
NOR2XL inst_cellmath__203_0_I2598 (.Y(N9265), .A(N7570), .B(N8696));
NOR2XL inst_cellmath__203_0_I2599 (.Y(N10020), .A(N7570), .B(N9044));
NOR2XL inst_cellmath__203_0_I2600 (.Y(N9035), .A(N7570), .B(N9436));
NOR2XL inst_cellmath__203_0_I2601 (.Y(N9810), .A(N7570), .B(N9816));
NOR2XL inst_cellmath__203_0_I2602 (.Y(N8827), .A(N7570), .B(N10177));
NOR2XL inst_cellmath__203_0_I2603 (.Y(N9592), .A(N7570), .B(N8837));
NOR2XL inst_cellmath__203_0_I2604 (.Y(N8642), .A(N7570), .B(N9206));
NOR2XL inst_cellmath__203_0_I2605 (.Y(N9359), .A(N7570), .B(N9598));
NOR2XL inst_cellmath__203_0_I2606 (.Y(N10104), .A(N7570), .B(N9967));
NOR2XL inst_cellmath__203_0_I2607 (.Y(N9131), .A(N7570), .B(N8646));
NOR2XL inst_cellmath__203_0_I2608 (.Y(N9898), .A(N7570), .B(N8985));
NOR2XL inst_cellmath__203_0_I2609 (.Y(N8915), .A(N7570), .B(N9366));
NOR2XL inst_cellmath__203_0_I2610 (.Y(N9683), .A(N7570), .B(N9753));
NOR2XL inst_cellmath__203_0_I2611 (.Y(N8714), .A(N7570), .B(N10112));
NOR2XL inst_cellmath__203_0_I2612 (.Y(N9835), .A(N7570), .B(N8772));
NOR2XL inst_cellmath__203_0_I2613 (.Y(N10193), .A(N7570), .B(N9136));
NOR2XL inst_cellmath__203_0_I2614 (.Y(N9226), .A(N7570), .B(N9527));
NOR2XL inst_cellmath__203_0_I2615 (.Y(N8784), .A(N7570), .B(N9907));
NOR2XL inst_cellmath__203_0_I2616 (.Y(N8754), .A(N7570), .B(N8595));
NOR2XL inst_cellmath__203_0_I2617 (.Y(N9775), .A(N7570), .B(N8923));
NAND2BX1 inst_cellmath__203_0_I2619 (.Y(N9073), .AN(inst_cellmath__61[2]), .B(inst_cellmath__61[1]));
NOR2XL inst_cellmath__203_0_I2621 (.Y(N8616), .A(N9664), .B(N7904));
MXI2XL inst_cellmath__203_0_I2622 (.Y(N10067), .A(N7390), .B(N9073), .S0(N8616));
MXI2XL inst_cellmath__203_0_I2623 (.Y(N10227), .A(N10030), .B(N9664), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2624 (.Y(N8734), .A(N7390), .B(N9073), .S0(N10227));
MXI2XL inst_cellmath__203_0_I2625 (.Y(N10167), .A(N8696), .B(N10030), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2626 (.Y(N9094), .A(N7390), .B(N9073), .S0(N10167));
MXI2XL inst_cellmath__203_0_I2627 (.Y(N10105), .A(N9044), .B(N8696), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2628 (.Y(N9485), .A(N7390), .B(N9073), .S0(N10105));
MXI2XL inst_cellmath__203_0_I2629 (.Y(N10045), .A(N9436), .B(N9044), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2630 (.Y(N9863), .A(N7390), .B(N9073), .S0(N10045));
MXI2XL inst_cellmath__203_0_I2631 (.Y(N9984), .A(N9816), .B(N9436), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2632 (.Y(N10218), .A(N7390), .B(N9073), .S0(N9984));
MXI2XL inst_cellmath__203_0_I2633 (.Y(N9924), .A(N10177), .B(N9816), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2634 (.Y(N8876), .A(N7390), .B(N9073), .S0(N9924));
MXI2XL inst_cellmath__203_0_I2635 (.Y(N9864), .A(N8837), .B(N10177), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2636 (.Y(N9258), .A(N7390), .B(N9073), .S0(N9864));
MXI2XL inst_cellmath__203_0_I2637 (.Y(N9802), .A(N9206), .B(N8837), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2638 (.Y(N9647), .A(N7390), .B(N9073), .S0(N9802));
MXI2XL inst_cellmath__203_0_I2639 (.Y(N9738), .A(N9598), .B(N9206), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2640 (.Y(N10009), .A(N7390), .B(N9073), .S0(N9738));
MXI2XL inst_cellmath__203_0_I2641 (.Y(N9677), .A(N9967), .B(N9598), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2642 (.Y(N8680), .A(N7390), .B(N9073), .S0(N9677));
MXI2XL inst_cellmath__203_0_I2643 (.Y(N9610), .A(N8646), .B(N9967), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2644 (.Y(N9028), .A(N7390), .B(N9073), .S0(N9610));
MXI2XL inst_cellmath__203_0_I2645 (.Y(N9542), .A(N8985), .B(N8646), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2646 (.Y(N9417), .A(N7390), .B(N9073), .S0(N9542));
MXI2XL inst_cellmath__203_0_I2647 (.Y(N9478), .A(N9366), .B(N8985), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2648 (.Y(N9801), .A(N7390), .B(N9073), .S0(N9478));
MXI2XL inst_cellmath__203_0_I2649 (.Y(N9410), .A(N9753), .B(N9366), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2650 (.Y(N10161), .A(N7390), .B(N9073), .S0(N9410));
MXI2XL inst_cellmath__203_0_I2651 (.Y(N9344), .A(N10112), .B(N9753), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2652 (.Y(N8818), .A(N7390), .B(N9073), .S0(N9344));
MXI2XL inst_cellmath__203_0_I2653 (.Y(N9278), .A(N8772), .B(N10112), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2654 (.Y(N9190), .A(N7390), .B(N9073), .S0(N9278));
MXI2XL inst_cellmath__203_0_I2655 (.Y(N9210), .A(N9136), .B(N8772), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2656 (.Y(N9582), .A(N7390), .B(N9073), .S0(N9210));
MXI2XL inst_cellmath__203_0_I2657 (.Y(N9144), .A(N9527), .B(N9136), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2658 (.Y(N9947), .A(N7390), .B(N9073), .S0(N9144));
MXI2XL inst_cellmath__203_0_I2659 (.Y(N9079), .A(N9907), .B(N9527), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2660 (.Y(N8632), .A(N7390), .B(N9073), .S0(N9079));
MXI2XL inst_cellmath__203_0_I2661 (.Y(N9016), .A(N8595), .B(N9907), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2662 (.Y(N8970), .A(N7390), .B(N9073), .S0(N9016));
MXI2XL inst_cellmath__203_0_I2663 (.Y(N8956), .A(N8923), .B(N8595), .S0(N7904));
MXI2XL inst_cellmath__203_0_I2664 (.Y(N9350), .A(N7390), .B(N9073), .S0(N8956));
NOR2BX1 inst_cellmath__203_0_I2665 (.Y(N8892), .AN(N7904), .B(N8923));
MXI2XL inst_cellmath__203_0_I2666 (.Y(N9736), .A(N7390), .B(N9073), .S0(N8892));
XNOR2X1 inst_cellmath__203_0_I2667 (.Y(N9514), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
NOR2XL inst_cellmath__203_0_I2668 (.Y(N9596), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
OAI2BB1X1 inst_cellmath__203_0_I2669 (.Y(N9124), .A0N(inst_cellmath__61[3]), .A1N(inst_cellmath__61[2]), .B0(inst_cellmath__61[4]));
INVXL inst_cellmath__203_0_I2670 (.Y(N9846), .A(N9124));
OR2XL inst_cellmath__203_0_I2671 (.Y(N9235), .A(N9596), .B(inst_cellmath__61[4]));
INVXL inst_cellmath__203_0_I2672 (.Y(N9626), .A(N9846));
NOR2XL inst_cellmath__203_0_I2673 (.Y(N8593), .A(N9664), .B(N9514));
MXI2XL inst_cellmath__203_0_I2674 (.Y(N10041), .A(N9626), .B(N9235), .S0(N8593));
MXI2XL inst_cellmath__203_0_I2675 (.Y(N10199), .A(N10030), .B(N9664), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2676 (.Y(N8707), .A(N9626), .B(N9235), .S0(N10199));
MXI2XL inst_cellmath__203_0_I2677 (.Y(N10138), .A(N8696), .B(N10030), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2678 (.Y(N9059), .A(N9626), .B(N9235), .S0(N10138));
MXI2XL inst_cellmath__203_0_I2679 (.Y(N10074), .A(N9044), .B(N8696), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2680 (.Y(N9450), .A(N9626), .B(N9235), .S0(N10074));
MXI2XL inst_cellmath__203_0_I2681 (.Y(N10019), .A(N9436), .B(N9044), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2682 (.Y(N9825), .A(N9626), .B(N9235), .S0(N10019));
MXI2XL inst_cellmath__203_0_I2683 (.Y(N9957), .A(N9816), .B(N9436), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2684 (.Y(N10187), .A(N9626), .B(N9235), .S0(N9957));
MXI2XL inst_cellmath__203_0_I2685 (.Y(N9897), .A(N10177), .B(N9816), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2686 (.Y(N8847), .A(N9626), .B(N9235), .S0(N9897));
MXI2XL inst_cellmath__203_0_I2687 (.Y(N9834), .A(N8837), .B(N10177), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2688 (.Y(N9216), .A(N9626), .B(N9235), .S0(N9834));
MXI2XL inst_cellmath__203_0_I2689 (.Y(N9773), .A(N9206), .B(N8837), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2690 (.Y(N9609), .A(N9626), .B(N9235), .S0(N9773));
MXI2XL inst_cellmath__203_0_I2691 (.Y(N9708), .A(N9598), .B(N9206), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2692 (.Y(N9977), .A(N9626), .B(N9235), .S0(N9708));
MXI2XL inst_cellmath__203_0_I2693 (.Y(N9645), .A(N9967), .B(N9598), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2694 (.Y(N8657), .A(N9626), .B(N9235), .S0(N9645));
MXI2XL inst_cellmath__203_0_I2695 (.Y(N9579), .A(N8646), .B(N9967), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2696 (.Y(N8998), .A(N9626), .B(N9235), .S0(N9579));
MXI2XL inst_cellmath__203_0_I2697 (.Y(N9511), .A(N8985), .B(N8646), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2698 (.Y(N9380), .A(N9626), .B(N9235), .S0(N9511));
MXI2XL inst_cellmath__203_0_I2699 (.Y(N9448), .A(N9366), .B(N8985), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2700 (.Y(N9764), .A(N9626), .B(N9235), .S0(N9448));
MXI2XL inst_cellmath__203_0_I2701 (.Y(N9378), .A(N9753), .B(N9366), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2702 (.Y(N10124), .A(N9626), .B(N9235), .S0(N9378));
MXI2XL inst_cellmath__203_0_I2703 (.Y(N9313), .A(N10112), .B(N9753), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2704 (.Y(N8785), .A(N9626), .B(N9235), .S0(N9313));
MXI2XL inst_cellmath__203_0_I2705 (.Y(N9249), .A(N8772), .B(N10112), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2706 (.Y(N9151), .A(N9626), .B(N9235), .S0(N9249));
MXI2XL inst_cellmath__203_0_I2707 (.Y(N9179), .A(N9136), .B(N8772), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2708 (.Y(N9541), .A(N9626), .B(N9235), .S0(N9179));
MXI2XL inst_cellmath__203_0_I2709 (.Y(N9112), .A(N9527), .B(N9136), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2710 (.Y(N9915), .A(N9626), .B(N9235), .S0(N9112));
MXI2XL inst_cellmath__203_0_I2711 (.Y(N9048), .A(N9907), .B(N9527), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2712 (.Y(N8603), .A(N9626), .B(N9235), .S0(N9048));
MXI2XL inst_cellmath__203_0_I2713 (.Y(N8988), .A(N8595), .B(N9907), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2714 (.Y(N8937), .A(N9626), .B(N9235), .S0(N8988));
MXI2XL inst_cellmath__203_0_I2715 (.Y(N8927), .A(N8923), .B(N8595), .S0(N9514));
MXI2XL inst_cellmath__203_0_I2716 (.Y(N9315), .A(N9626), .B(N9235), .S0(N8927));
NOR2BX1 inst_cellmath__203_0_I2717 (.Y(N8864), .AN(N9514), .B(N8923));
MXI2XL inst_cellmath__203_0_I2718 (.Y(N9702), .A(N9626), .B(N9235), .S0(N8864));
XNOR2X1 inst_cellmath__203_0_I2719 (.Y(N9477), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
NOR2XL inst_cellmath__203_0_I2720 (.Y(N9562), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
OAI2BB1X1 inst_cellmath__203_0_I2721 (.Y(N9086), .A0N(inst_cellmath__61[5]), .A1N(inst_cellmath__61[4]), .B0(inst_cellmath__61[6]));
INVXL inst_cellmath__203_0_I2722 (.Y(N9993), .A(N9086));
OR2XL inst_cellmath__203_0_I2723 (.Y(N9396), .A(N9562), .B(inst_cellmath__61[6]));
INVXL inst_cellmath__203_0_I2724 (.Y(N9785), .A(N9993));
NOR2XL inst_cellmath__203_0_I2725 (.Y(N10229), .A(N9664), .B(N9477));
MXI2XL inst_cellmath__203_0_I2726 (.Y(N10003), .A(N9785), .B(N9396), .S0(N10229));
MXI2XL inst_cellmath__203_0_I2727 (.Y(N10171), .A(N10030), .B(N9664), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2728 (.Y(N8676), .A(N9785), .B(N9396), .S0(N10171));
MXI2XL inst_cellmath__203_0_I2729 (.Y(N10107), .A(N8696), .B(N10030), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2730 (.Y(N9023), .A(N9785), .B(N9396), .S0(N10107));
MXI2XL inst_cellmath__203_0_I2731 (.Y(N10048), .A(N9044), .B(N8696), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2732 (.Y(N9408), .A(N9785), .B(N9396), .S0(N10048));
MXI2XL inst_cellmath__203_0_I2733 (.Y(N9986), .A(N9436), .B(N9044), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2734 (.Y(N9793), .A(N9785), .B(N9396), .S0(N9986));
MXI2XL inst_cellmath__203_0_I2735 (.Y(N9927), .A(N9816), .B(N9436), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2736 (.Y(N10153), .A(N9785), .B(N9396), .S0(N9927));
MXI2XL inst_cellmath__203_0_I2737 (.Y(N9868), .A(N10177), .B(N9816), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2738 (.Y(N8812), .A(N9785), .B(N9396), .S0(N9868));
MXI2XL inst_cellmath__203_0_I2739 (.Y(N9804), .A(N8837), .B(N10177), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2740 (.Y(N9181), .A(N9785), .B(N9396), .S0(N9804));
MXI2XL inst_cellmath__203_0_I2741 (.Y(N9741), .A(N9206), .B(N8837), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2742 (.Y(N9572), .A(N9785), .B(N9396), .S0(N9741));
MXI2XL inst_cellmath__203_0_I2743 (.Y(N9680), .A(N9598), .B(N9206), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2744 (.Y(N9941), .A(N9785), .B(N9396), .S0(N9680));
MXI2XL inst_cellmath__203_0_I2745 (.Y(N9612), .A(N9967), .B(N9598), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2746 (.Y(N8626), .A(N9785), .B(N9396), .S0(N9612));
MXI2XL inst_cellmath__203_0_I2747 (.Y(N9545), .A(N8646), .B(N9967), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2748 (.Y(N8962), .A(N9785), .B(N9396), .S0(N9545));
MXI2XL inst_cellmath__203_0_I2749 (.Y(N9482), .A(N8985), .B(N8646), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2750 (.Y(N9342), .A(N9785), .B(N9396), .S0(N9482));
MXI2XL inst_cellmath__203_0_I2751 (.Y(N9413), .A(N9366), .B(N8985), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2752 (.Y(N9728), .A(N9785), .B(N9396), .S0(N9413));
MXI2XL inst_cellmath__203_0_I2753 (.Y(N9347), .A(N9753), .B(N9366), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2754 (.Y(N10090), .A(N9785), .B(N9396), .S0(N9347));
MXI2XL inst_cellmath__203_0_I2755 (.Y(N9282), .A(N10112), .B(N9753), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2756 (.Y(N8753), .A(N9785), .B(N9396), .S0(N9282));
MXI2XL inst_cellmath__203_0_I2757 (.Y(N9212), .A(N8772), .B(N10112), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2758 (.Y(N9114), .A(N9785), .B(N9396), .S0(N9212));
MXI2XL inst_cellmath__203_0_I2759 (.Y(N9146), .A(N9136), .B(N8772), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2760 (.Y(N9504), .A(N9785), .B(N9396), .S0(N9146));
MXI2XL inst_cellmath__203_0_I2761 (.Y(N9081), .A(N9527), .B(N9136), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2762 (.Y(N9884), .A(N9785), .B(N9396), .S0(N9081));
MXI2XL inst_cellmath__203_0_I2763 (.Y(N9018), .A(N9907), .B(N9527), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2764 (.Y(N10237), .A(N9785), .B(N9396), .S0(N9018));
MXI2XL inst_cellmath__203_0_I2765 (.Y(N8958), .A(N8595), .B(N9907), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2766 (.Y(N8901), .A(N9785), .B(N9396), .S0(N8958));
MXI2XL inst_cellmath__203_0_I2767 (.Y(N8894), .A(N8923), .B(N8595), .S0(N9477));
MXI2XL inst_cellmath__203_0_I2768 (.Y(N9276), .A(N9785), .B(N9396), .S0(N8894));
NOR2BX1 inst_cellmath__203_0_I2769 (.Y(N8836), .AN(N9477), .B(N8923));
MXI2XL inst_cellmath__203_0_I2770 (.Y(N9668), .A(N9785), .B(N9396), .S0(N8836));
XNOR2X1 inst_cellmath__203_0_I2771 (.Y(N9441), .A(inst_cellmath__61[7]), .B(inst_cellmath__61[6]));
NOR2XL inst_cellmath__203_0_I2772 (.Y(N9528), .A(inst_cellmath__61[7]), .B(inst_cellmath__61[6]));
OAI2BB1X1 inst_cellmath__203_0_I2773 (.Y(N9050), .A0N(inst_cellmath__61[7]), .A1N(inst_cellmath__61[6]), .B0(inst_cellmath__61[8]));
INVXL inst_cellmath__203_0_I2774 (.Y(N10142), .A(N9050));
OR2XL inst_cellmath__203_0_I2775 (.Y(N9560), .A(N9528), .B(inst_cellmath__61[8]));
INVXL inst_cellmath__203_0_I2776 (.Y(N9932), .A(N10142));
NOR2XL inst_cellmath__203_0_I2777 (.Y(N10202), .A(N9664), .B(N9441));
MXI2XL inst_cellmath__203_0_I2778 (.Y(N9970), .A(N9932), .B(N9560), .S0(N10202));
MXI2XL inst_cellmath__203_0_I2779 (.Y(N10141), .A(N10030), .B(N9664), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2780 (.Y(N8650), .A(N9932), .B(N9560), .S0(N10141));
MXI2XL inst_cellmath__203_0_I2781 (.Y(N10076), .A(N8696), .B(N10030), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2782 (.Y(N8990), .A(N9932), .B(N9560), .S0(N10076));
MXI2XL inst_cellmath__203_0_I2783 (.Y(N10022), .A(N9044), .B(N8696), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2784 (.Y(N9371), .A(N9932), .B(N9560), .S0(N10022));
MXI2XL inst_cellmath__203_0_I2785 (.Y(N9959), .A(N9436), .B(N9044), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2786 (.Y(N9756), .A(N9932), .B(N9560), .S0(N9959));
MXI2XL inst_cellmath__203_0_I2787 (.Y(N9900), .A(N9816), .B(N9436), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2788 (.Y(N10118), .A(N9932), .B(N9560), .S0(N9900));
MXI2XL inst_cellmath__203_0_I2789 (.Y(N9836), .A(N10177), .B(N9816), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2790 (.Y(N8778), .A(N9932), .B(N9560), .S0(N9836));
MXI2XL inst_cellmath__203_0_I2791 (.Y(N9776), .A(N8837), .B(N10177), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2792 (.Y(N9141), .A(N9932), .B(N9560), .S0(N9776));
MXI2XL inst_cellmath__203_0_I2793 (.Y(N9710), .A(N9206), .B(N8837), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2794 (.Y(N9533), .A(N9932), .B(N9560), .S0(N9710));
MXI2XL inst_cellmath__203_0_I2795 (.Y(N9648), .A(N9598), .B(N9206), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2796 (.Y(N9910), .A(N9932), .B(N9560), .S0(N9648));
MXI2XL inst_cellmath__203_0_I2797 (.Y(N9583), .A(N9967), .B(N9598), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2798 (.Y(N8597), .A(N9932), .B(N9560), .S0(N9583));
MXI2XL inst_cellmath__203_0_I2799 (.Y(N9515), .A(N8646), .B(N9967), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2800 (.Y(N8928), .A(N9932), .B(N9560), .S0(N9515));
MXI2XL inst_cellmath__203_0_I2801 (.Y(N9451), .A(N8985), .B(N8646), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2802 (.Y(N9306), .A(N9932), .B(N9560), .S0(N9451));
MXI2XL inst_cellmath__203_0_I2803 (.Y(N9381), .A(N9366), .B(N8985), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2804 (.Y(N9693), .A(N9932), .B(N9560), .S0(N9381));
MXI2XL inst_cellmath__203_0_I2805 (.Y(N9316), .A(N9753), .B(N9366), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2806 (.Y(N10058), .A(N9932), .B(N9560), .S0(N9316));
MXI2XL inst_cellmath__203_0_I2807 (.Y(N9251), .A(N10112), .B(N9753), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2808 (.Y(N8723), .A(N9932), .B(N9560), .S0(N9251));
MXI2XL inst_cellmath__203_0_I2809 (.Y(N9182), .A(N8772), .B(N10112), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2810 (.Y(N9077), .A(N9932), .B(N9560), .S0(N9182));
MXI2XL inst_cellmath__203_0_I2811 (.Y(N9115), .A(N9136), .B(N8772), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2812 (.Y(N9470), .A(N9932), .B(N9560), .S0(N9115));
MXI2XL inst_cellmath__203_0_I2813 (.Y(N9051), .A(N9527), .B(N9136), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2814 (.Y(N9851), .A(N9932), .B(N9560), .S0(N9051));
MXI2XL inst_cellmath__203_0_I2815 (.Y(N8991), .A(N9907), .B(N9527), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2816 (.Y(N10206), .A(N9932), .B(N9560), .S0(N8991));
MXI2XL inst_cellmath__203_0_I2817 (.Y(N8929), .A(N8595), .B(N9907), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2818 (.Y(N8866), .A(N9932), .B(N9560), .S0(N8929));
MXI2XL inst_cellmath__203_0_I2819 (.Y(N8867), .A(N8923), .B(N8595), .S0(N9441));
MXI2XL inst_cellmath__203_0_I2820 (.Y(N9242), .A(N9932), .B(N9560), .S0(N8867));
NOR2BX1 inst_cellmath__203_0_I2821 (.Y(N8805), .AN(N9441), .B(N8923));
MXI2XL inst_cellmath__203_0_I2822 (.Y(N9630), .A(N9932), .B(N9560), .S0(N8805));
XNOR2X1 inst_cellmath__203_0_I2823 (.Y(N9399), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
NOR2XL inst_cellmath__203_0_I2824 (.Y(N9497), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
OAI2BB1X1 inst_cellmath__203_0_I2825 (.Y(N9013), .A0N(inst_cellmath__61[9]), .A1N(inst_cellmath__61[8]), .B0(inst_cellmath__61[10]));
INVXL inst_cellmath__203_0_I2826 (.Y(N8617), .A(N9013));
OR2XL inst_cellmath__203_0_I2827 (.Y(N9718), .A(N9497), .B(inst_cellmath__61[10]));
INVXL inst_cellmath__203_0_I2828 (.Y(N10077), .A(N8617));
NOR2XL inst_cellmath__203_0_I2829 (.Y(N10175), .A(N9664), .B(N9399));
MXI2XL inst_cellmath__203_0_I2830 (.Y(N9936), .A(N10077), .B(N9718), .S0(N10175));
MXI2XL inst_cellmath__203_0_I2831 (.Y(N10110), .A(N10030), .B(N9664), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2832 (.Y(N8620), .A(N10077), .B(N9718), .S0(N10110));
MXI2XL inst_cellmath__203_0_I2833 (.Y(N10052), .A(N8696), .B(N10030), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2834 (.Y(N8955), .A(N10077), .B(N9718), .S0(N10052));
MXI2XL inst_cellmath__203_0_I2835 (.Y(N9990), .A(N9044), .B(N8696), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2836 (.Y(N9333), .A(N10077), .B(N9718), .S0(N9990));
MXI2XL inst_cellmath__203_0_I2837 (.Y(N9929), .A(N9436), .B(N9044), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2838 (.Y(N9721), .A(N10077), .B(N9718), .S0(N9929));
MXI2XL inst_cellmath__203_0_I2839 (.Y(N9872), .A(N9816), .B(N9436), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2840 (.Y(N10083), .A(N10077), .B(N9718), .S0(N9872));
MXI2XL inst_cellmath__203_0_I2841 (.Y(N9808), .A(N10177), .B(N9816), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2842 (.Y(N8744), .A(N10077), .B(N9718), .S0(N9808));
MXI2XL inst_cellmath__203_0_I2843 (.Y(N9745), .A(N8837), .B(N10177), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2844 (.Y(N9104), .A(N10077), .B(N9718), .S0(N9745));
MXI2XL inst_cellmath__203_0_I2845 (.Y(N9682), .A(N9206), .B(N8837), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2846 (.Y(N9496), .A(N10077), .B(N9718), .S0(N9682));
MXI2XL inst_cellmath__203_0_I2847 (.Y(N9616), .A(N9598), .B(N9206), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2848 (.Y(N9877), .A(N10077), .B(N9718), .S0(N9616));
MXI2XL inst_cellmath__203_0_I2849 (.Y(N9549), .A(N9967), .B(N9598), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2850 (.Y(N10230), .A(N10077), .B(N9718), .S0(N9549));
MXI2XL inst_cellmath__203_0_I2851 (.Y(N9484), .A(N8646), .B(N9967), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2852 (.Y(N8891), .A(N10077), .B(N9718), .S0(N9484));
MXI2XL inst_cellmath__203_0_I2853 (.Y(N9416), .A(N8985), .B(N8646), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2854 (.Y(N9267), .A(N10077), .B(N9718), .S0(N9416));
MXI2XL inst_cellmath__203_0_I2855 (.Y(N9349), .A(N9366), .B(N8985), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2856 (.Y(N9661), .A(N10077), .B(N9718), .S0(N9349));
MXI2XL inst_cellmath__203_0_I2857 (.Y(N9284), .A(N9753), .B(N9366), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2858 (.Y(N10027), .A(N10077), .B(N9718), .S0(N9284));
MXI2XL inst_cellmath__203_0_I2859 (.Y(N9215), .A(N10112), .B(N9753), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2860 (.Y(N8692), .A(N10077), .B(N9718), .S0(N9215));
MXI2XL inst_cellmath__203_0_I2861 (.Y(N9150), .A(N8772), .B(N10112), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2862 (.Y(N9040), .A(N10077), .B(N9718), .S0(N9150));
MXI2XL inst_cellmath__203_0_I2863 (.Y(N9084), .A(N9136), .B(N8772), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2864 (.Y(N9432), .A(N10077), .B(N9718), .S0(N9084));
MXI2XL inst_cellmath__203_0_I2865 (.Y(N9020), .A(N9527), .B(N9136), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2866 (.Y(N9813), .A(N10077), .B(N9718), .S0(N9020));
MXI2XL inst_cellmath__203_0_I2867 (.Y(N8961), .A(N9907), .B(N9527), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2868 (.Y(N10173), .A(N10077), .B(N9718), .S0(N8961));
MXI2XL inst_cellmath__203_0_I2869 (.Y(N8899), .A(N8595), .B(N9907), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2870 (.Y(N8834), .A(N10077), .B(N9718), .S0(N8899));
MXI2XL inst_cellmath__203_0_I2871 (.Y(N8840), .A(N8923), .B(N8595), .S0(N9399));
MXI2XL inst_cellmath__203_0_I2872 (.Y(N9200), .A(N10077), .B(N9718), .S0(N8840));
NOR2BX1 inst_cellmath__203_0_I2873 (.Y(N8776), .AN(N9399), .B(N8923));
MXI2XL inst_cellmath__203_0_I2874 (.Y(N9595), .A(N10077), .B(N9718), .S0(N8776));
XNOR2X1 inst_cellmath__203_0_I2875 (.Y(N9364), .A(inst_cellmath__61[11]), .B(inst_cellmath__61[10]));
NOR2XL inst_cellmath__203_0_I2876 (.Y(N9468), .A(inst_cellmath__61[11]), .B(inst_cellmath__61[10]));
OAI2BB1X1 inst_cellmath__203_0_I2877 (.Y(N8982), .A0N(inst_cellmath__61[11]), .A1N(inst_cellmath__61[10]), .B0(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I2878 (.Y(N8742), .A(N8982));
OR2XL inst_cellmath__203_0_I2879 (.Y(N9874), .A(N9468), .B(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I2880 (.Y(N10228), .A(N8742));
NOR2XL inst_cellmath__203_0_I2881 (.Y(N10146), .A(N9664), .B(N9364));
MXI2XL inst_cellmath__203_0_I2882 (.Y(N9904), .A(N10228), .B(N9874), .S0(N10146));
MXI2XL inst_cellmath__203_0_I2883 (.Y(N10080), .A(N10030), .B(N9664), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2884 (.Y(N8591), .A(N10228), .B(N9874), .S0(N10080));
MXI2XL inst_cellmath__203_0_I2885 (.Y(N10025), .A(N8696), .B(N10030), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2886 (.Y(N8919), .A(N10228), .B(N9874), .S0(N10025));
MXI2XL inst_cellmath__203_0_I2887 (.Y(N9962), .A(N9044), .B(N8696), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2888 (.Y(N9297), .A(N10228), .B(N9874), .S0(N9962));
MXI2XL inst_cellmath__203_0_I2889 (.Y(N9902), .A(N9436), .B(N9044), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2890 (.Y(N9686), .A(N10228), .B(N9874), .S0(N9902));
MXI2XL inst_cellmath__203_0_I2891 (.Y(N9839), .A(N9816), .B(N9436), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2892 (.Y(N10050), .A(N10228), .B(N9874), .S0(N9839));
MXI2XL inst_cellmath__203_0_I2893 (.Y(N9778), .A(N10177), .B(N9816), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2894 (.Y(N8717), .A(N10228), .B(N9874), .S0(N9778));
MXI2XL inst_cellmath__203_0_I2895 (.Y(N9714), .A(N8837), .B(N10177), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2896 (.Y(N9067), .A(N10228), .B(N9874), .S0(N9714));
MXI2XL inst_cellmath__203_0_I2897 (.Y(N9652), .A(N9206), .B(N8837), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2898 (.Y(N9460), .A(N10228), .B(N9874), .S0(N9652));
MXI2XL inst_cellmath__203_0_I2899 (.Y(N9586), .A(N9598), .B(N9206), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2900 (.Y(N9842), .A(N10228), .B(N9874), .S0(N9586));
MXI2XL inst_cellmath__203_0_I2901 (.Y(N9518), .A(N9967), .B(N9598), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2902 (.Y(N10197), .A(N10228), .B(N9874), .S0(N9518));
MXI2XL inst_cellmath__203_0_I2903 (.Y(N9454), .A(N8646), .B(N9967), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2904 (.Y(N8857), .A(N10228), .B(N9874), .S0(N9454));
MXI2XL inst_cellmath__203_0_I2905 (.Y(N9384), .A(N8985), .B(N8646), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2906 (.Y(N9231), .A(N10228), .B(N9874), .S0(N9384));
MXI2XL inst_cellmath__203_0_I2907 (.Y(N9319), .A(N9366), .B(N8985), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2908 (.Y(N9621), .A(N10228), .B(N9874), .S0(N9319));
MXI2XL inst_cellmath__203_0_I2909 (.Y(N9254), .A(N9753), .B(N9366), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2910 (.Y(N9988), .A(N10228), .B(N9874), .S0(N9254));
MXI2XL inst_cellmath__203_0_I2911 (.Y(N9185), .A(N10112), .B(N9753), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2912 (.Y(N8668), .A(N10228), .B(N9874), .S0(N9185));
MXI2XL inst_cellmath__203_0_I2913 (.Y(N9118), .A(N8772), .B(N10112), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2914 (.Y(N9005), .A(N10228), .B(N9874), .S0(N9118));
MXI2XL inst_cellmath__203_0_I2915 (.Y(N9055), .A(N9136), .B(N8772), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2916 (.Y(N9392), .A(N10228), .B(N9874), .S0(N9055));
MXI2XL inst_cellmath__203_0_I2917 (.Y(N8995), .A(N9527), .B(N9136), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2918 (.Y(N9781), .A(N10228), .B(N9874), .S0(N8995));
MXI2XL inst_cellmath__203_0_I2919 (.Y(N8932), .A(N9907), .B(N9527), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2920 (.Y(N10135), .A(N10228), .B(N9874), .S0(N8932));
MXI2XL inst_cellmath__203_0_I2921 (.Y(N8869), .A(N8595), .B(N9907), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2922 (.Y(N8797), .A(N10228), .B(N9874), .S0(N8869));
MXI2XL inst_cellmath__203_0_I2923 (.Y(N8807), .A(N8923), .B(N8595), .S0(N9364));
MXI2XL inst_cellmath__203_0_I2924 (.Y(N9166), .A(N10228), .B(N9874), .S0(N8807));
NOR2BX1 inst_cellmath__203_0_I2925 (.Y(N8748), .AN(N9364), .B(N8923));
MXI2XL inst_cellmath__203_0_I2926 (.Y(N9555), .A(N10228), .B(N9874), .S0(N8748));
XNOR2X1 inst_cellmath__203_0_I2927 (.Y(N9330), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
NOR2XL inst_cellmath__203_0_I2928 (.Y(N9435), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
OAI2BB1X1 inst_cellmath__203_0_I2929 (.Y(N8946), .A0N(inst_cellmath__61[13]), .A1N(inst_cellmath__61[12]), .B0(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I2930 (.Y(N8886), .A(N8946));
OR2XL inst_cellmath__203_0_I2931 (.Y(N10023), .A(N9435), .B(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I2932 (.Y(N8689), .A(N8886));
NOR2XL inst_cellmath__203_0_I2933 (.Y(N10113), .A(N9664), .B(N9330));
MXI2XL inst_cellmath__203_0_I2934 (.Y(N9870), .A(N8689), .B(N10023), .S0(N10113));
MXI2XL inst_cellmath__203_0_I2935 (.Y(N10054), .A(N10030), .B(N9664), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2936 (.Y(N10224), .A(N8689), .B(N10023), .S0(N10054));
MXI2XL inst_cellmath__203_0_I2937 (.Y(N9994), .A(N8696), .B(N10030), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2938 (.Y(N8881), .A(N8689), .B(N10023), .S0(N9994));
MXI2XL inst_cellmath__203_0_I2939 (.Y(N9933), .A(N9044), .B(N8696), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2940 (.Y(N9262), .A(N8689), .B(N10023), .S0(N9933));
MXI2XL inst_cellmath__203_0_I2941 (.Y(N9875), .A(N9436), .B(N9044), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2942 (.Y(N9655), .A(N8689), .B(N10023), .S0(N9875));
MXI2XL inst_cellmath__203_0_I2943 (.Y(N9811), .A(N9816), .B(N9436), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2944 (.Y(N10016), .A(N8689), .B(N10023), .S0(N9811));
MXI2XL inst_cellmath__203_0_I2945 (.Y(N9747), .A(N10177), .B(N9816), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2946 (.Y(N8686), .A(N8689), .B(N10023), .S0(N9747));
MXI2XL inst_cellmath__203_0_I2947 (.Y(N9684), .A(N8837), .B(N10177), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2948 (.Y(N9031), .A(N8689), .B(N10023), .S0(N9684));
MXI2XL inst_cellmath__203_0_I2949 (.Y(N9618), .A(N9206), .B(N8837), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2950 (.Y(N9422), .A(N8689), .B(N10023), .S0(N9618));
MXI2XL inst_cellmath__203_0_I2951 (.Y(N9552), .A(N9598), .B(N9206), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2952 (.Y(N9806), .A(N8689), .B(N10023), .S0(N9552));
MXI2XL inst_cellmath__203_0_I2953 (.Y(N9487), .A(N9967), .B(N9598), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2954 (.Y(N10164), .A(N8689), .B(N10023), .S0(N9487));
MXI2XL inst_cellmath__203_0_I2955 (.Y(N9419), .A(N8646), .B(N9967), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2956 (.Y(N8826), .A(N8689), .B(N10023), .S0(N9419));
MXI2XL inst_cellmath__203_0_I2957 (.Y(N9353), .A(N8985), .B(N8646), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2958 (.Y(N9195), .A(N8689), .B(N10023), .S0(N9353));
MXI2XL inst_cellmath__203_0_I2959 (.Y(N9286), .A(N9366), .B(N8985), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2960 (.Y(N9588), .A(N8689), .B(N10023), .S0(N9286));
MXI2XL inst_cellmath__203_0_I2961 (.Y(N9218), .A(N9753), .B(N9366), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2962 (.Y(N9956), .A(N8689), .B(N10023), .S0(N9218));
MXI2XL inst_cellmath__203_0_I2963 (.Y(N9153), .A(N10112), .B(N9753), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2964 (.Y(N8638), .A(N8689), .B(N10023), .S0(N9153));
MXI2XL inst_cellmath__203_0_I2965 (.Y(N9087), .A(N8772), .B(N10112), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2966 (.Y(N8974), .A(N8689), .B(N10023), .S0(N9087));
MXI2XL inst_cellmath__203_0_I2967 (.Y(N9024), .A(N9136), .B(N8772), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2968 (.Y(N9358), .A(N8689), .B(N10023), .S0(N9024));
MXI2XL inst_cellmath__203_0_I2969 (.Y(N8963), .A(N9527), .B(N9136), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2970 (.Y(N9742), .A(N8689), .B(N10023), .S0(N8963));
MXI2XL inst_cellmath__203_0_I2971 (.Y(N8902), .A(N9907), .B(N9527), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2972 (.Y(N10100), .A(N8689), .B(N10023), .S0(N8902));
MXI2XL inst_cellmath__203_0_I2973 (.Y(N8842), .A(N8595), .B(N9907), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2974 (.Y(N8766), .A(N8689), .B(N10023), .S0(N8842));
MXI2XL inst_cellmath__203_0_I2975 (.Y(N8779), .A(N8923), .B(N8595), .S0(N9330));
MXI2XL inst_cellmath__203_0_I2976 (.Y(N9128), .A(N8689), .B(N10023), .S0(N8779));
NOR2BX1 inst_cellmath__203_0_I2977 (.Y(N8724), .AN(N9330), .B(N8923));
MXI2XL inst_cellmath__203_0_I2978 (.Y(N9628), .A(N8689), .B(N10023), .S0(N8724));
XNOR2X1 inst_cellmath__203_0_I2979 (.Y(N9290), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
NOR2XL inst_cellmath__203_0_I2980 (.Y(N9401), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
OAI2BB1X1 inst_cellmath__203_0_I2981 (.Y(N8912), .A0N(inst_cellmath__61[15]), .A1N(inst_cellmath__61[14]), .B0(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I2982 (.Y(N9036), .A(N8912));
OR2XL inst_cellmath__203_0_I2983 (.Y(N10168), .A(N9401), .B(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I2984 (.Y(inst_cellmath__203__W0[42]), .A(N9036));
NOR2XL inst_cellmath__203_0_I2985 (.Y(N10084), .A(N9664), .B(N9290));
MXI2XL inst_cellmath__203_0_I2986 (.Y(N9833), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N10084));
MXI2XL inst_cellmath__203_0_I2987 (.Y(N10028), .A(N10030), .B(N9664), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2988 (.Y(N10190), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N10028));
MXI2XL inst_cellmath__203_0_I2989 (.Y(N9965), .A(N8696), .B(N10030), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2990 (.Y(N8850), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9965));
MXI2XL inst_cellmath__203_0_I2991 (.Y(N9905), .A(N9044), .B(N8696), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2992 (.Y(N9224), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9905));
MXI2XL inst_cellmath__203_0_I2993 (.Y(N9843), .A(N9436), .B(N9044), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2994 (.Y(N9613), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9843));
MXI2XL inst_cellmath__203_0_I2995 (.Y(N9782), .A(N9816), .B(N9436), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2996 (.Y(N9980), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9782));
MXI2XL inst_cellmath__203_0_I2997 (.Y(N9716), .A(N10177), .B(N9816), .S0(N9290));
MXI2XL inst_cellmath__203_0_I2998 (.Y(N8662), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9716));
MXI2XL inst_cellmath__203_0_I2999 (.Y(N9656), .A(N8837), .B(N10177), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3000 (.Y(N9000), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9656));
MXI2XL inst_cellmath__203_0_I3001 (.Y(N9590), .A(N9206), .B(N8837), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3002 (.Y(N9386), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9590));
MXI2XL inst_cellmath__203_0_I3003 (.Y(N9520), .A(N9598), .B(N9206), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3004 (.Y(N9772), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9520));
MXI2XL inst_cellmath__203_0_I3005 (.Y(N9457), .A(N9967), .B(N9598), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3006 (.Y(N10128), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9457));
MXI2XL inst_cellmath__203_0_I3007 (.Y(N9388), .A(N8646), .B(N9967), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3008 (.Y(N8789), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9388));
MXI2XL inst_cellmath__203_0_I3009 (.Y(N9323), .A(N8985), .B(N8646), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3010 (.Y(N9158), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9323));
MXI2XL inst_cellmath__203_0_I3011 (.Y(N9256), .A(N9366), .B(N8985), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3012 (.Y(N9546), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9256));
MXI2XL inst_cellmath__203_0_I3013 (.Y(N9188), .A(N9753), .B(N9366), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3014 (.Y(N9920), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9188));
MXI2XL inst_cellmath__203_0_I3015 (.Y(N9122), .A(N10112), .B(N9753), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3016 (.Y(N8609), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9122));
MXI2XL inst_cellmath__203_0_I3017 (.Y(N9057), .A(N8772), .B(N10112), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3018 (.Y(N8940), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N9057));
MXI2XL inst_cellmath__203_0_I3019 (.Y(N8997), .A(N9136), .B(N8772), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3020 (.Y(N9321), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8997));
MXI2XL inst_cellmath__203_0_I3021 (.Y(N8935), .A(N9527), .B(N9136), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3022 (.Y(N9707), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8935));
MXI2XL inst_cellmath__203_0_I3023 (.Y(N8871), .A(N9907), .B(N9527), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3024 (.Y(N10066), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8871));
MXI2XL inst_cellmath__203_0_I3025 (.Y(N8811), .A(N8595), .B(N9907), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3026 (.Y(N8732), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8811));
MXI2XL inst_cellmath__203_0_I3027 (.Y(N8752), .A(N8923), .B(N8595), .S0(N9290));
MXI2XL inst_cellmath__203_0_I3028 (.Y(N9092), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8752));
NOR2BX1 inst_cellmath__203_0_I3029 (.Y(N8700), .AN(N9290), .B(N8923));
MXI2XL inst_cellmath__203_0_I3030 (.Y(inst_cellmath__203__W1[42]), .A(inst_cellmath__203__W0[42]), .B(N10168), .S0(N8700));
ADDHX1 inst_cellmath__203_0_I3031 (.CO(inst_cellmath__203__W0[2]), .S(inst_cellmath__203__W1[1]), .A(N10207), .B(inst_cellmath__198[19]));
ADDHX1 inst_cellmath__203_0_I3032 (.CO(inst_cellmath__203__W0[3]), .S(inst_cellmath__203__W1[2]), .A(N9240), .B(N9295));
ADDHX1 inst_cellmath__203_0_I3033 (.CO(N10211), .S(N9855), .A(N9998), .B(N9696));
ADDFX1 inst_cellmath__203_0_I3034 (.CO(inst_cellmath__203__W0[4]), .S(inst_cellmath__203__W1[3]), .A(N9871), .B(N9687), .CI(N9855));
ADDFX1 inst_cellmath__203_0_I3035 (.CO(N10001), .S(N9638), .A(N9014), .B(N9492), .CI(N10051));
ADDFX1 inst_cellmath__203_0_I3036 (.CO(inst_cellmath__203__W0[5]), .S(inst_cellmath__203__W1[4]), .A(N10211), .B(N10222), .CI(N9638));
ADDFX1 inst_cellmath__203_0_I3037 (.CO(N9791), .S(N9405), .A(N10226), .B(inst_cellmath__61[2]), .CI(N10067));
ADDFX1 inst_cellmath__203_0_I3038 (.CO(N8808), .S(N10151), .A(N9787), .B(N9405), .CI(N8716));
ADDFX1 inst_cellmath__203_0_I3039 (.CO(N9570), .S(N9177), .A(N8882), .B(N9853), .CI(N9062));
ADDFX1 inst_cellmath__203_0_I3040 (.CO(inst_cellmath__203__W0[6]), .S(inst_cellmath__203__W1[5]), .A(N10151), .B(N10001), .CI(N9177));
ADDFX1 inst_cellmath__203_0_I3041 (.CO(N9339), .S(N8960), .A(N8734), .B(N9265), .CI(N9791));
ADDFX1 inst_cellmath__203_0_I3042 (.CO(N10089), .S(N9725), .A(N8804), .B(N8960), .CI(N9068));
ADDFX1 inst_cellmath__203_0_I3043 (.CO(N9110), .S(N8749), .A(N9456), .B(N9263), .CI(N8808));
ADDFX1 inst_cellmath__203_0_I3044 (.CO(inst_cellmath__203__W0[7]), .S(inst_cellmath__203__W1[6]), .A(N9570), .B(N9725), .CI(N8749));
ADDFX1 inst_cellmath__203_0_I3045 (.CO(N8898), .S(N10234), .A(N10020), .B(N9846), .CI(N10041));
ADDFX1 inst_cellmath__203_0_I3046 (.CO(N9665), .S(N9273), .A(N10234), .B(N9094), .CI(N9339));
ADDFX1 inst_cellmath__203_0_I3047 (.CO(N8697), .S(N10033), .A(N9563), .B(N9273), .CI(N9461));
ADDFX1 inst_cellmath__203_0_I3048 (.CO(N9439), .S(N9046), .A(N9653), .B(N10000), .CI(N9831));
ADDFX1 inst_cellmath__203_0_I3049 (.CO(N10179), .S(N9817), .A(N10089), .B(N10007), .CI(N10033));
ADDFX1 inst_cellmath__203_0_I3050 (.CO(inst_cellmath__203__W0[8]), .S(inst_cellmath__203__W1[7]), .A(N9046), .B(N9110), .CI(N9817));
ADDFX1 inst_cellmath__203_0_I3051 (.CO(N9968), .S(N9599), .A(N8707), .B(N9035), .CI(N9485));
ADDFX1 inst_cellmath__203_0_I3052 (.CO(N8987), .S(N8647), .A(N9599), .B(N8898), .CI(N9665));
ADDFX1 inst_cellmath__203_0_I3053 (.CO(N9754), .S(N9369), .A(N8621), .B(N8647), .CI(N9840));
ADDFX1 inst_cellmath__203_0_I3054 (.CO(N8775), .S(N10115), .A(N10191), .B(N10017), .CI(N8679));
ADDFX1 inst_cellmath__203_0_I3055 (.CO(N9530), .S(N9137), .A(N9369), .B(N8697), .CI(N9439));
ADDFX1 inst_cellmath__203_0_I3056 (.CO(inst_cellmath__203__W0[9]), .S(inst_cellmath__203__W1[8]), .A(N10115), .B(N10179), .CI(N9137));
ADDFX1 inst_cellmath__203_0_I3057 (.CO(N9303), .S(N8925), .A(N9810), .B(N9993), .CI(N10003));
ADDFX1 inst_cellmath__203_0_I3058 (.CO(N10056), .S(N9692), .A(N9863), .B(N9059), .CI(N9968));
ADDFX1 inst_cellmath__203_0_I3059 (.CO(N9076), .S(N8721), .A(N9692), .B(N8925), .CI(N8987));
ADDFX1 inst_cellmath__203_0_I3060 (.CO(N9848), .S(N9465), .A(N8721), .B(N9334), .CI(N10148));
ADDFX1 inst_cellmath__203_0_I3061 (.CO(N8862), .S(N10204), .A(N9214), .B(N10198), .CI(N8687));
ADDFX1 inst_cellmath__203_0_I3062 (.CO(N9629), .S(N9237), .A(N9026), .B(N8851), .CI(N9754));
ADDFX1 inst_cellmath__203_0_I3063 (.CO(N8671), .S(N9995), .A(N8775), .B(N9465), .CI(N10204));
ADDFX1 inst_cellmath__203_0_I3064 (.CO(inst_cellmath__203__W0[10]), .S(inst_cellmath__203__W1[9]), .A(N9530), .B(N9237), .CI(N9995));
ADDFX1 inst_cellmath__203_0_I3065 (.CO(N10144), .S(N9786), .A(N8676), .B(N8827), .CI(N9450));
ADDFX1 inst_cellmath__203_0_I3066 (.CO(N9171), .S(N8802), .A(N9303), .B(N10218), .CI(N9786));
ADDFX1 inst_cellmath__203_0_I3067 (.CO(N9934), .S(N9561), .A(N8802), .B(N10056), .CI(N9076));
ADDFX1 inst_cellmath__203_0_I3068 (.CO(N8952), .S(N8618), .A(N9561), .B(N10081), .CI(N8858));
ADDFX1 inst_cellmath__203_0_I3069 (.CO(N9719), .S(N9332), .A(N9032), .B(N9606), .CI(N9222));
ADDFX1 inst_cellmath__203_0_I3070 (.CO(N8743), .S(N10079), .A(N9848), .B(N9414), .CI(N8618));
ADDFX1 inst_cellmath__203_0_I3071 (.CO(N9494), .S(N9100), .A(N9629), .B(N8862), .CI(N9332));
ADDFX1 inst_cellmath__203_0_I3072 (.CO(inst_cellmath__203__W0[11]), .S(inst_cellmath__203__W1[10]), .A(N8671), .B(N10079), .CI(N9100));
ADDFX1 inst_cellmath__203_0_I3073 (.CO(N9266), .S(N8888), .A(N9592), .B(N10142), .CI(N9970));
ADDFX1 inst_cellmath__203_0_I3074 (.CO(N10024), .S(N9658), .A(N9825), .B(N9023), .CI(N8876));
ADDFX1 inst_cellmath__203_0_I3075 (.CO(N9037), .S(N8690), .A(N8888), .B(N10144), .CI(N9658));
ADDFX1 inst_cellmath__203_0_I3076 (.CO(N9812), .S(N9428), .A(N8690), .B(N9171), .CI(N9105));
ADDFX1 inst_cellmath__203_0_I3077 (.CO(N8831), .S(N10169), .A(N9428), .B(N9934), .CI(N9229));
ADDFX1 inst_cellmath__203_0_I3078 (.CO(N9593), .S(N9198), .A(N9975), .B(N8623), .CI(N9423));
ADDFX1 inst_cellmath__203_0_I3079 (.CO(N8643), .S(N9961), .A(N10149), .B(N9614), .CI(N9798));
ADDFX1 inst_cellmath__203_0_I3080 (.CO(N9361), .S(N8978), .A(N10169), .B(N8952), .CI(N9719));
ADDFX1 inst_cellmath__203_0_I3081 (.CO(N10106), .S(N9748), .A(N8743), .B(N9198), .CI(N9961));
ADDFX1 inst_cellmath__203_0_I3082 (.CO(inst_cellmath__203__W0[12]), .S(inst_cellmath__203__W1[11]), .A(N9494), .B(N8978), .CI(N9748));
ADDFX1 inst_cellmath__203_0_I3083 (.CO(N9901), .S(N9522), .A(N8650), .B(N8642), .CI(N9408));
ADDFX1 inst_cellmath__203_0_I3084 (.CO(N8916), .S(N8589), .A(N9258), .B(N10187), .CI(N9266));
ADDFX1 inst_cellmath__203_0_I3085 (.CO(N9685), .S(N9293), .A(N9522), .B(N10024), .CI(N8589));
ADDFX1 inst_cellmath__203_0_I3086 (.CO(N8715), .S(N10046), .A(N9293), .B(N9037), .CI(N9878));
ADDFX1 inst_cellmath__203_0_I3087 (.CO(N9458), .S(N9065), .A(N10046), .B(N9812), .CI(N9622));
ADDFX1 inst_cellmath__203_0_I3088 (.CO(N10195), .S(N9838), .A(N9807), .B(N8655), .CI(N9981));
ADDFX1 inst_cellmath__203_0_I3089 (.CO(N9227), .S(N8854), .A(N8809), .B(N10156), .CI(N8831));
ADDFX1 inst_cellmath__203_0_I3090 (.CO(N9985), .S(N9619), .A(N9593), .B(N9065), .CI(N8643));
ADDFX1 inst_cellmath__203_0_I3091 (.CO(N9004), .S(N8665), .A(N8854), .B(N9838), .CI(N9361));
ADDFX1 inst_cellmath__203_0_I3092 (.CO(inst_cellmath__203__W0[13]), .S(inst_cellmath__203__W1[12]), .A(N10106), .B(N9619), .CI(N8665));
ADDFX1 inst_cellmath__203_0_I3093 (.CO(N8793), .S(N10132), .A(N9359), .B(N8617), .CI(N9936));
ADDFX1 inst_cellmath__203_0_I3094 (.CO(N9553), .S(N9162), .A(N9647), .B(N8990), .CI(N9793));
ADDFX1 inst_cellmath__203_0_I3095 (.CO(N8611), .S(N9925), .A(N9901), .B(N8847), .CI(N10132));
ADDFX1 inst_cellmath__203_0_I3096 (.CO(N9326), .S(N8945), .A(N9162), .B(N8916), .CI(N9925));
ADDFX1 inst_cellmath__203_0_I3097 (.CO(N10072), .S(N9712), .A(N8945), .B(N9685), .CI(N8890));
ADDFX1 inst_cellmath__203_0_I3098 (.CO(N9096), .S(N8736), .A(N9712), .B(N8715), .CI(N9989));
ADDFX1 inst_cellmath__203_0_I3099 (.CO(N9865), .S(N9490), .A(N8747), .B(N8996), .CI(N9178));
ADDFX1 inst_cellmath__203_0_I3100 (.CO(N8880), .S(N10220), .A(N8659), .B(N10165), .CI(N8816));
ADDFX1 inst_cellmath__203_0_I3101 (.CO(N9650), .S(N9259), .A(N9458), .B(N9367), .CI(N8736));
ADDFX1 inst_cellmath__203_0_I3102 (.CO(N8682), .S(N10014), .A(N9227), .B(N10195), .CI(N9490));
ADDFX1 inst_cellmath__203_0_I3103 (.CO(N9421), .S(N9030), .A(N9985), .B(N10220), .CI(N9259));
ADDFX1 inst_cellmath__203_0_I3104 (.CO(inst_cellmath__203__W0[14]), .S(inst_cellmath__203__W1[13]), .A(N10014), .B(N9004), .CI(N9030));
ADDFX1 inst_cellmath__203_0_I3105 (.CO(N9192), .S(N8822), .A(N8620), .B(N10104), .CI(N9371));
ADDFX1 inst_cellmath__203_0_I3106 (.CO(N9952), .S(N9585), .A(N10009), .B(N10153), .CI(N9216));
ADDFX1 inst_cellmath__203_0_I3107 (.CO(N8972), .S(N8635), .A(N9553), .B(N8793), .CI(N8822));
ADDFX1 inst_cellmath__203_0_I3108 (.CO(N9739), .S(N9355), .A(N8611), .B(N9585), .CI(N8635));
ADDFX1 inst_cellmath__203_0_I3109 (.CO(N8762), .S(N10098), .A(N9355), .B(N9326), .CI(N9662));
ADDFX1 inst_cellmath__203_0_I3110 (.CO(N9517), .S(N9126), .A(N10098), .B(N10072), .CI(N8666));
ADDFX1 inst_cellmath__203_0_I3111 (.CO(N8583), .S(N9893), .A(N8823), .B(N9377), .CI(N9001));
ADDFX1 inst_cellmath__203_0_I3112 (.CO(N9288), .S(N8910), .A(N9568), .B(N9187), .CI(N9755));
ADDFX1 inst_cellmath__203_0_I3113 (.CO(N10043), .S(N9678), .A(N9126), .B(N9096), .CI(N9865));
ADDFX1 inst_cellmath__203_0_I3114 (.CO(N9060), .S(N8710), .A(N9893), .B(N8880), .CI(N9650));
ADDFX1 inst_cellmath__203_0_I3115 (.CO(N9829), .S(N9453), .A(N9678), .B(N8910), .CI(N8682));
ADDFX1 inst_cellmath__203_0_I3116 (.CO(inst_cellmath__203__W0[15]), .S(inst_cellmath__203__W1[14]), .A(N9421), .B(N8710), .CI(N9453));
ADDHX1 inst_cellmath__203_0_I3117 (.CO(N9611), .S(N9221), .A(N8742), .B(N9131));
ADDFX1 inst_cellmath__203_0_I3118 (.CO(N8658), .S(N9978), .A(N9221), .B(N9904), .CI(N8955));
ADDFX1 inst_cellmath__203_0_I3119 (.CO(N9383), .S(N8999), .A(N9756), .B(N9609), .CI(N8812));
ADDFX1 inst_cellmath__203_0_I3120 (.CO(N10126), .S(N9768), .A(N9192), .B(N8680), .CI(N9952));
ADDFX1 inst_cellmath__203_0_I3121 (.CO(N9155), .S(N8787), .A(N8999), .B(N9978), .CI(N8972));
ADDFX1 inst_cellmath__203_0_I3122 (.CO(N9917), .S(N9543), .A(N8787), .B(N9768), .CI(N9739));
ADDFX1 inst_cellmath__203_0_I3123 (.CO(N8938), .S(N8605), .A(N9543), .B(N8693), .CI(N8762));
ADDFX1 inst_cellmath__203_0_I3124 (.CO(N9704), .S(N9318), .A(N10078), .B(N8605), .CI(N9006));
ADDFX1 inst_cellmath__203_0_I3125 (.CO(N8730), .S(N10064), .A(N9196), .B(N9761), .CI(N9387));
ADDFX1 inst_cellmath__203_0_I3126 (.CO(N9480), .S(N9089), .A(N9939), .B(N9577), .CI(N10116));
ADDFX1 inst_cellmath__203_0_I3127 (.CO(N10214), .S(N9859), .A(N9318), .B(N9517), .CI(N8583));
ADDFX1 inst_cellmath__203_0_I3128 (.CO(N9253), .S(N8873), .A(N10064), .B(N9288), .CI(N9089));
ADDFX1 inst_cellmath__203_0_I3129 (.CO(N10005), .S(N9642), .A(N9859), .B(N10043), .CI(N9060));
ADDFX1 inst_cellmath__203_0_I3130 (.CO(inst_cellmath__203__W0[16]), .S(inst_cellmath__203__W1[15]), .A(N8873), .B(N9829), .CI(N9642));
ADDFX1 inst_cellmath__203_0_I3131 (.CO(N9794), .S(N9411), .A(N9611), .B(N9898), .CI(N8591));
ADDFX1 inst_cellmath__203_0_I3132 (.CO(N8814), .S(N10155), .A(N10118), .B(N9333), .CI(N9181));
ADDFX1 inst_cellmath__203_0_I3133 (.CO(N9575), .S(N9183), .A(N9028), .B(N9977), .CI(N8658));
ADDFX1 inst_cellmath__203_0_I3134 (.CO(N8627), .S(N9944), .A(N9411), .B(N9383), .CI(N10155));
ADDFX1 inst_cellmath__203_0_I3135 (.CO(N9346), .S(N8965), .A(N9183), .B(N10126), .CI(N9944));
ADDFX1 inst_cellmath__203_0_I3136 (.CO(N10092), .S(N9730), .A(N9430), .B(N9155), .CI(N8965));
ADDFX1 inst_cellmath__203_0_I3137 (.CO(N9116), .S(N8756), .A(N9730), .B(N9917), .CI(N8938));
ADDFX1 inst_cellmath__203_0_I3138 (.CO(N9887), .S(N9507), .A(N8756), .B(N9101), .CI(N9393));
ADDFX1 inst_cellmath__203_0_I3139 (.CO(N8904), .S(N10238), .A(N9589), .B(N10122), .CI(N9770));
ADDFX1 inst_cellmath__203_0_I3140 (.CO(N9670), .S(N9280), .A(N8625), .B(N9945), .CI(N8773));
ADDFX1 inst_cellmath__203_0_I3141 (.CO(N8703), .S(N10035), .A(N9507), .B(N9704), .CI(N8730));
ADDFX1 inst_cellmath__203_0_I3142 (.CO(N9443), .S(N9052), .A(N10238), .B(N9480), .CI(N9280));
ADDFX1 inst_cellmath__203_0_I3143 (.CO(N10182), .S(N9821), .A(N10035), .B(N10214), .CI(N9253));
ADDFX1 inst_cellmath__203_0_I3144 (.CO(inst_cellmath__203__W0[17]), .S(inst_cellmath__203__W1[16]), .A(N10005), .B(N9052), .CI(N9821));
ADDFX1 inst_cellmath__203_0_I3145 (.CO(N9971), .S(N9602), .A(N8915), .B(N8886), .CI(N9870));
ADDFX1 inst_cellmath__203_0_I3146 (.CO(N8992), .S(N8653), .A(N9572), .B(N9417), .CI(N8919));
ADDFX1 inst_cellmath__203_0_I3147 (.CO(N9759), .S(N9373), .A(N8778), .B(N9721), .CI(N8657));
ADDFX1 inst_cellmath__203_0_I3148 (.CO(N8780), .S(N10119), .A(N8814), .B(N9794), .CI(N9602));
ADDFX1 inst_cellmath__203_0_I3149 (.CO(N9535), .S(N9145), .A(N9575), .B(N8653), .CI(N9373));
ADDFX1 inst_cellmath__203_0_I3150 (.CO(N8598), .S(N9911), .A(N10119), .B(N8627), .CI(N9145));
ADDFX1 inst_cellmath__203_0_I3151 (.CO(N9308), .S(N8930), .A(N10174), .B(N9346), .CI(N9911));
ADDFX1 inst_cellmath__203_0_I3152 (.CO(N10059), .S(N9695), .A(N8930), .B(N10092), .CI(N9116));
ADDFX1 inst_cellmath__203_0_I3153 (.CO(N9080), .S(N8725), .A(N9779), .B(N9876), .CI(N8783));
ADDFX1 inst_cellmath__203_0_I3154 (.CO(N9852), .S(N9472), .A(N9695), .B(N9954), .CI(N8959));
ADDFX1 inst_cellmath__203_0_I3155 (.CO(N8868), .S(N10209), .A(N8630), .B(N10129), .CI(N9138));
ADDFX1 inst_cellmath__203_0_I3156 (.CO(N9633), .S(N9244), .A(N8904), .B(N9887), .CI(N8725));
ADDFX1 inst_cellmath__203_0_I3157 (.CO(N8673), .S(N9999), .A(N9472), .B(N9670), .CI(N10209));
ADDFX1 inst_cellmath__203_0_I3158 (.CO(N9402), .S(N9017), .A(N9244), .B(N8703), .CI(N9443));
ADDFX1 inst_cellmath__203_0_I3159 (.CO(inst_cellmath__203__W0[18]), .S(inst_cellmath__203__W1[17]), .A(N10182), .B(N9999), .CI(N9017));
ADDFX1 inst_cellmath__203_0_I3160 (.CO(N9175), .S(N8806), .A(N10224), .B(N9683), .CI(N9297));
ADDFX1 inst_cellmath__203_0_I3161 (.CO(N9937), .S(N9566), .A(N10083), .B(N9801), .CI(N9141));
ADDFX1 inst_cellmath__203_0_I3162 (.CO(N8957), .S(N8622), .A(N8998), .B(N9941), .CI(N9971));
ADDFX1 inst_cellmath__203_0_I3163 (.CO(N9722), .S(N9337), .A(N9759), .B(N8992), .CI(N8806));
ADDFX1 inst_cellmath__203_0_I3164 (.CO(N8746), .S(N10085), .A(N8622), .B(N9566), .CI(N8780));
ADDFX1 inst_cellmath__203_0_I3165 (.CO(N9499), .S(N9107), .A(N9337), .B(N9535), .CI(N10085));
ADDFX1 inst_cellmath__203_0_I3166 (.CO(N10231), .S(N9880), .A(N9201), .B(N8598), .CI(N9107));
ADDFX1 inst_cellmath__203_0_I3167 (.CO(N9270), .S(N8893), .A(N9880), .B(N9308), .CI(N8887));
ADDFX1 inst_cellmath__203_0_I3168 (.CO(N10029), .S(N9663), .A(N10136), .B(N10059), .CI(N9148));
ADDFX1 inst_cellmath__203_0_I3169 (.CO(N9042), .S(N8695), .A(N8790), .B(N8639), .CI(N9340));
ADDFX1 inst_cellmath__203_0_I3170 (.CO(N9815), .S(N9434), .A(N8893), .B(N8966), .CI(N9531));
ADDFX1 inst_cellmath__203_0_I3171 (.CO(N8835), .S(N10176), .A(N9852), .B(N9080), .CI(N9663));
ADDFX1 inst_cellmath__203_0_I3172 (.CO(N9597), .S(N9205), .A(N8695), .B(N8868), .CI(N9434));
ADDFX1 inst_cellmath__203_0_I3173 (.CO(N8645), .S(N9966), .A(N10176), .B(N9633), .CI(N8673));
ADDFX1 inst_cellmath__203_0_I3174 (.CO(inst_cellmath__203__W0[19]), .S(inst_cellmath__203__W1[18]), .A(N9402), .B(N9205), .CI(N9966));
ADDFX1 inst_cellmath__203_0_I3175 (.CO(N10111), .S(N9752), .A(N8714), .B(N9036), .CI(N9833));
ADDFX1 inst_cellmath__203_0_I3176 (.CO(N9135), .S(N8771), .A(N9533), .B(N9380), .CI(N8881));
ADDFX1 inst_cellmath__203_0_I3177 (.CO(N9906), .S(N9526), .A(N9686), .B(N10161), .CI(N8744));
ADDFX1 inst_cellmath__203_0_I3178 (.CO(N8921), .S(N8594), .A(N9175), .B(N8626), .CI(N9937));
ADDFX1 inst_cellmath__203_0_I3179 (.CO(N9689), .S(N9299), .A(N8957), .B(N9752), .CI(N8771));
ADDFX1 inst_cellmath__203_0_I3180 (.CO(N8719), .S(N10053), .A(N9722), .B(N9526), .CI(N8594));
ADDFX1 inst_cellmath__203_0_I3181 (.CO(N9462), .S(N9072), .A(N8746), .B(N9299), .CI(N10053));
ADDFX1 inst_cellmath__203_0_I3182 (.CO(N10201), .S(N9845), .A(N9499), .B(N9963), .CI(N9072));
ADDFX1 inst_cellmath__203_0_I3183 (.CO(N9234), .S(N8860), .A(N9845), .B(N10231), .CI(N9659));
ADDFX1 inst_cellmath__203_0_I3184 (.CO(N9991), .S(N9625), .A(N9270), .B(N8798), .CI(N9537));
ADDFX1 inst_cellmath__203_0_I3185 (.CO(N9011), .S(N8670), .A(N9156), .B(N8975), .CI(N9726));
ADDFX1 inst_cellmath__203_0_I3186 (.CO(N9784), .S(N9394), .A(N8860), .B(N9348), .CI(N9908));
ADDFX1 inst_cellmath__203_0_I3187 (.CO(N8800), .S(N10140), .A(N9042), .B(N10029), .CI(N9625));
ADDFX1 inst_cellmath__203_0_I3188 (.CO(N9559), .S(N9169), .A(N8670), .B(N9815), .CI(N9394));
ADDFX1 inst_cellmath__203_0_I3189 (.CO(N8615), .S(N9930), .A(N10140), .B(N8835), .CI(N9597));
ADDFX1 inst_cellmath__203_0_I3190 (.CO(inst_cellmath__203__W0[20]), .S(inst_cellmath__203__W1[19]), .A(N8645), .B(N9169), .CI(N9930));
INVXL inst_cellmath__203_0_I3191 (.Y(N8649), .A(N9835));
ADDFX1 inst_cellmath__203_0_I3192 (.CO(N10075), .S(N9717), .A(N9262), .B(N10190), .CI(N8649));
ADDFX1 inst_cellmath__203_0_I3193 (.CO(N9873), .S(N9493), .A(N8818), .B(N9764), .CI(N10050));
ADDFX1 inst_cellmath__203_0_I3194 (.CO(N8885), .S(N10225), .A(N9104), .B(N9910), .CI(N8962));
ADDFX1 inst_cellmath__203_0_I3195 (.CO(N9657), .S(N9264), .A(N9135), .B(N10111), .CI(N9906));
ADDFX1 inst_cellmath__203_0_I3196 (.CO(N8688), .S(N10021), .A(N9493), .B(N9717), .CI(N10225));
ADDFX1 inst_cellmath__203_0_I3197 (.CO(N9426), .S(N9034), .A(N9689), .B(N8921), .CI(N9264));
ADDFX1 inst_cellmath__203_0_I3198 (.CO(N10166), .S(N9809), .A(N8719), .B(N10021), .CI(N9034));
ADDFX1 inst_cellmath__203_0_I3199 (.CO(N9197), .S(N8829), .A(N9462), .B(N9147), .CI(N9809));
ADDFX1 inst_cellmath__203_0_I3200 (.CO(N9958), .S(N9591), .A(N8829), .B(N10201), .CI(N8691));
ADDFX1 inst_cellmath__203_0_I3201 (.CO(N8977), .S(N8641), .A(N9234), .B(N9164), .CI(N9913));
ADDFX1 inst_cellmath__203_0_I3202 (.CO(N9746), .S(N9360), .A(N9547), .B(N9356), .CI(N10087));
ADDFX1 inst_cellmath__203_0_I3203 (.CO(N8768), .S(N10103), .A(N9591), .B(N9733), .CI(N8596));
ADDFX1 inst_cellmath__203_0_I3204 (.CO(N9521), .S(N9130), .A(N9011), .B(N9991), .CI(N8641));
ADDFX1 inst_cellmath__203_0_I3205 (.CO(N8588), .S(N9899), .A(N9360), .B(N9784), .CI(N10103));
ADDFX1 inst_cellmath__203_0_I3206 (.CO(N9291), .S(N8914), .A(N9130), .B(N8800), .CI(N9559));
ADDFX1 inst_cellmath__203_0_I3207 (.CO(inst_cellmath__203__W0[21]), .S(inst_cellmath__203__W1[20]), .A(N8615), .B(N9899), .CI(N8914));
ADDFX1 inst_cellmath__203_0_I3208 (.CO(N9064), .S(N8713), .A(N9190), .B(N10193), .CI(N8649));
ADDFX1 inst_cellmath__203_0_I3209 (.CO(N8852), .S(N10194), .A(N9496), .B(N9342), .CI(N8850));
ADDFX1 inst_cellmath__203_0_I3210 (.CO(N9617), .S(N9225), .A(N9655), .B(N10124), .CI(N8717));
ADDFX1 inst_cellmath__203_0_I3211 (.CO(N8663), .S(N9983), .A(N10075), .B(N8597), .CI(N9873));
ADDFX1 inst_cellmath__203_0_I3212 (.CO(N9389), .S(N9003), .A(N8713), .B(N8885), .CI(N10194));
ADDFX1 inst_cellmath__203_0_I3213 (.CO(N10131), .S(N9774), .A(N9657), .B(N9225), .CI(N9983));
ADDFX1 inst_cellmath__203_0_I3214 (.CO(N9159), .S(N8791), .A(N9003), .B(N8688), .CI(N9426));
ADDFX1 inst_cellmath__203_0_I3215 (.CO(N9923), .S(N9551), .A(N10166), .B(N9774), .CI(N8791));
ADDFX1 inst_cellmath__203_0_I3216 (.CO(N8943), .S(N8610), .A(N9551), .B(N9197), .CI(N9427));
ADDFX1 inst_cellmath__203_0_I3217 (.CO(N9709), .S(N9324), .A(N9958), .B(N9556), .CI(N8600));
ADDFX1 inst_cellmath__203_0_I3218 (.CO(N8733), .S(N10068), .A(N9921), .B(N9743), .CI(N8750));
ADDFX1 inst_cellmath__203_0_I3219 (.CO(N9486), .S(N9093), .A(N8610), .B(N10093), .CI(N8926));
ADDFX1 inst_cellmath__203_0_I3220 (.CO(N10217), .S(N9862), .A(N9746), .B(N8977), .CI(N9324));
ADDFX1 inst_cellmath__203_0_I3221 (.CO(N9257), .S(N8877), .A(N10068), .B(N8768), .CI(N9093));
ADDFX1 inst_cellmath__203_0_I3222 (.CO(N10011), .S(N9646), .A(N9862), .B(N9521), .CI(N8588));
ADDFX1 inst_cellmath__203_0_I3223 (.CO(inst_cellmath__203__W0[22]), .S(inst_cellmath__203__W1[21]), .A(N9291), .B(N8877), .CI(N9646));
ADDFX1 inst_cellmath__203_0_I3224 (.CO(N9800), .S(N9418), .A(N9226), .B(N9835), .CI(N9728));
ADDFX1 inst_cellmath__203_0_I3225 (.CO(N8820), .S(N10160), .A(N9224), .B(N8785), .CI(N10016));
ADDFX1 inst_cellmath__203_0_I3226 (.CO(N9581), .S(N9189), .A(N9067), .B(N9877), .CI(N8928));
ADDFX1 inst_cellmath__203_0_I3227 (.CO(N8631), .S(N9950), .A(N9064), .B(N9582), .CI(N8852));
ADDFX1 inst_cellmath__203_0_I3228 (.CO(N9352), .S(N8969), .A(N9418), .B(N9617), .CI(N10160));
ADDFX1 inst_cellmath__203_0_I3229 (.CO(N10096), .S(N9735), .A(N8663), .B(N9189), .CI(N9950));
ADDFX1 inst_cellmath__203_0_I3230 (.CO(N9123), .S(N8760), .A(N8969), .B(N9389), .CI(N10131));
ADDFX1 inst_cellmath__203_0_I3231 (.CO(N9891), .S(N9513), .A(N9159), .B(N9735), .CI(N8760));
ADDFX1 inst_cellmath__203_0_I3232 (.CO(N8908), .S(N8581), .A(N9513), .B(N9923), .CI(N8931));
ADDFX1 inst_cellmath__203_0_I3233 (.CO(N9676), .S(N9285), .A(N8943), .B(N10170), .CI(N8581));
ADDFX1 inst_cellmath__203_0_I3234 (.CO(N8708), .S(N10040), .A(N10101), .B(N8933), .CI(N8606));
ADDFX1 inst_cellmath__203_0_I3235 (.CO(N9449), .S(N9058), .A(N9111), .B(N8757), .CI(N9304));
ADDFX1 inst_cellmath__203_0_I3236 (.CO(N10186), .S(N9827), .A(N9285), .B(N9709), .CI(N8733));
ADDFX1 inst_cellmath__203_0_I3237 (.CO(N9217), .S(N8846), .A(N10040), .B(N9486), .CI(N9058));
ADDFX1 inst_cellmath__203_0_I3238 (.CO(N9976), .S(N9608), .A(N9827), .B(N10217), .CI(N9257));
ADDFX1 inst_cellmath__203_0_I3239 (.CO(inst_cellmath__203__W0[23]), .S(inst_cellmath__203__W1[22]), .A(N10011), .B(N8846), .CI(N9608));
INVXL inst_cellmath__203_0_I3240 (.Y(N10205), .A(N8784));
ADDFX1 inst_cellmath__203_0_I3241 (.CO(N9766), .S(N9379), .A(N9306), .B(N9151), .CI(N10205));
ADDFX1 inst_cellmath__203_0_I3242 (.CO(N9540), .S(N9152), .A(N9460), .B(N10090), .CI(N9613));
ADDFX1 inst_cellmath__203_0_I3243 (.CO(N8602), .S(N9914), .A(N8686), .B(N9947), .CI(N10230));
ADDFX1 inst_cellmath__203_0_I3244 (.CO(N9314), .S(N8936), .A(N8820), .B(N9800), .CI(N9581));
ADDFX1 inst_cellmath__203_0_I3245 (.CO(N10063), .S(N9701), .A(N9152), .B(N9379), .CI(N9914));
ADDFX1 inst_cellmath__203_0_I3246 (.CO(N9085), .S(N8728), .A(N9352), .B(N8631), .CI(N8936));
ADDFX1 inst_cellmath__203_0_I3247 (.CO(N9857), .S(N9479), .A(N10096), .B(N9701), .CI(N8728));
ADDFX1 inst_cellmath__203_0_I3248 (.CO(N8872), .S(N10212), .A(N9479), .B(N9123), .CI(N9891));
ADDFX1 inst_cellmath__203_0_I3249 (.CO(N9639), .S(N9250), .A(N9199), .B(N10212), .CI(N8908));
ADDFX1 inst_cellmath__203_0_I3250 (.CO(N8675), .S(N10004), .A(N8763), .B(N9312), .CI(N8941));
ADDFX1 inst_cellmath__203_0_I3251 (.CO(N9409), .S(N9022), .A(N9500), .B(N9120), .CI(N9690));
ADDFX1 inst_cellmath__203_0_I3252 (.CO(N10152), .S(N9792), .A(N9676), .B(N9250), .CI(N8708));
ADDFX1 inst_cellmath__203_0_I3253 (.CO(N9180), .S(N8813), .A(N10004), .B(N9449), .CI(N9022));
ADDFX1 inst_cellmath__203_0_I3254 (.CO(N9942), .S(N9571), .A(N9792), .B(N10186), .CI(N9217));
ADDFX1 inst_cellmath__203_0_I3255 (.CO(inst_cellmath__203__W0[24]), .S(inst_cellmath__203__W1[23]), .A(N9976), .B(N8813), .CI(N9571));
INVXL inst_cellmath__203_0_I3256 (.Y(N10145), .A(N8754));
ADDFX1 inst_cellmath__203_0_I3257 (.CO(N9727), .S(N9343), .A(N9693), .B(N8784), .CI(N10145));
ADDFX1 inst_cellmath__203_0_I3258 (.CO(N9503), .S(N9113), .A(N9980), .B(N8753), .CI(N9541));
ADDFX1 inst_cellmath__203_0_I3259 (.CO(N10236), .S(N9885), .A(N9842), .B(N8632), .CI(N9031));
ADDFX1 inst_cellmath__203_0_I3260 (.CO(N9277), .S(N8900), .A(N9766), .B(N8891), .CI(N9540));
ADDFX1 inst_cellmath__203_0_I3261 (.CO(N10034), .S(N9667), .A(N9343), .B(N8602), .CI(N9113));
ADDFX1 inst_cellmath__203_0_I3262 (.CO(N9049), .S(N8701), .A(N9314), .B(N9885), .CI(N8900));
ADDFX1 inst_cellmath__203_0_I3263 (.CO(N9819), .S(N9440), .A(N9667), .B(N10063), .CI(N9085));
ADDFX1 inst_cellmath__203_0_I3264 (.CO(N8841), .S(N10181), .A(N9857), .B(N8701), .CI(N9440));
ADDFX1 inst_cellmath__203_0_I3265 (.CO(N9600), .S(N9209), .A(N8872), .B(N10181), .CI(N9082));
ADDFX1 inst_cellmath__203_0_I3266 (.CO(N8651), .S(N9969), .A(N9209), .B(N9960), .CI(N9697));
ADDFX1 inst_cellmath__203_0_I3267 (.CO(N9370), .S(N8989), .A(N9882), .B(N9639), .CI(N9509));
ADDFX1 inst_cellmath__203_0_I3268 (.CO(N10117), .S(N9757), .A(N10057), .B(N9322), .CI(N8675));
ADDFX1 inst_cellmath__203_0_I3269 (.CO(N9143), .S(N8777), .A(N9409), .B(N9969), .CI(N8989));
ADDFX1 inst_cellmath__203_0_I3270 (.CO(N9909), .S(N9532), .A(N9757), .B(N10152), .CI(N9180));
ADDFX1 inst_cellmath__203_0_I3271 (.CO(inst_cellmath__203__W0[25]), .S(inst_cellmath__203__W1[24]), .A(N9942), .B(N8777), .CI(N9532));
XNOR2X1 inst_cellmath__203_0_I3272 (.Y(N9305), .A(N9775), .B(N8754));
OR2XL inst_cellmath__203_0_I3273 (.Y(N9694), .A(N9775), .B(N8754));
ADDFX1 inst_cellmath__203_0_I3274 (.CO(N9469), .S(N9078), .A(N9114), .B(N9305), .CI(N9422));
ADDFX1 inst_cellmath__203_0_I3275 (.CO(N10208), .S(N9850), .A(N10058), .B(N9267), .CI(N8970));
ADDFX1 inst_cellmath__203_0_I3276 (.CO(N9241), .S(N8865), .A(N8662), .B(N9915), .CI(N10197));
ADDFX1 inst_cellmath__203_0_I3277 (.CO(N9997), .S(N9631), .A(N9503), .B(N9727), .CI(N10236));
ADDFX1 inst_cellmath__203_0_I3278 (.CO(N9015), .S(N8672), .A(N9850), .B(N9078), .CI(N8865));
ADDFX1 inst_cellmath__203_0_I3279 (.CO(N9788), .S(N9398), .A(N10034), .B(N9277), .CI(N9631));
ADDFX1 inst_cellmath__203_0_I3280 (.CO(N8803), .S(N10147), .A(N9049), .B(N8672), .CI(N9398));
ADDFX1 inst_cellmath__203_0_I3281 (.CO(N9564), .S(N9173), .A(N10147), .B(N9819), .CI(N8841));
ADDFX1 inst_cellmath__203_0_I3282 (.CO(N8619), .S(N9935), .A(N9173), .B(N8979), .CI(N9600));
ADDFX1 inst_cellmath__203_0_I3283 (.CO(N9336), .S(N8954), .A(N9706), .B(N10060), .CI(N10235));
ADDFX1 inst_cellmath__203_0_I3284 (.CO(N10082), .S(N9720), .A(N8722), .B(N9888), .CI(N9935));
ADDFX1 inst_cellmath__203_0_I3285 (.CO(N9103), .S(N8745), .A(N9370), .B(N8651), .CI(N8954));
ADDFX1 inst_cellmath__203_0_I3286 (.CO(N9879), .S(N9495), .A(N9720), .B(N10117), .CI(N9143));
ADDFX1 inst_cellmath__203_0_I3287 (.CO(inst_cellmath__203__W0[26]), .S(inst_cellmath__203__W1[25]), .A(N9909), .B(N8745), .CI(N9495));
ADDHX1 inst_cellmath__203_0_I3288 (.CO(N9660), .S(N9269), .A(N9694), .B(N9350));
ADDFX1 inst_cellmath__203_0_I3289 (.CO(N8694), .S(N10026), .A(N9661), .B(N9269), .CI(N8723));
ADDFX1 inst_cellmath__203_0_I3290 (.CO(N9431), .S(N9039), .A(N9806), .B(N8603), .CI(N9000));
ADDFX1 inst_cellmath__203_0_I3291 (.CO(N10172), .S(N9814), .A(N8857), .B(N9504), .CI(N9469));
ADDFX1 inst_cellmath__203_0_I3292 (.CO(N9203), .S(N8833), .A(N9241), .B(N10208), .CI(N10026));
ADDFX1 inst_cellmath__203_0_I3293 (.CO(N9964), .S(N9594), .A(N9997), .B(N9039), .CI(N9814));
ADDFX1 inst_cellmath__203_0_I3294 (.CO(N8981), .S(N8644), .A(N8833), .B(N9015), .CI(N9788));
ADDFX1 inst_cellmath__203_0_I3295 (.CO(N9751), .S(N9363), .A(N8644), .B(N9594), .CI(N8803));
ADDFX1 inst_cellmath__203_0_I3296 (.CO(N8770), .S(N10108), .A(N9564), .B(N9363), .CI(N9246));
ADDFX1 inst_cellmath__203_0_I3297 (.CO(N9525), .S(N9133), .A(N10108), .B(N9749), .CI(N8727));
ADDFX1 inst_cellmath__203_0_I3298 (.CO(N8592), .S(N9903), .A(N8896), .B(N8580), .CI(N8619));
ADDFX1 inst_cellmath__203_0_I3299 (.CO(N9296), .S(N8918), .A(N9336), .B(N9074), .CI(N9133));
ADDFX1 inst_cellmath__203_0_I3300 (.CO(N10049), .S(N9688), .A(N9903), .B(N10082), .CI(N9103));
ADDFX1 inst_cellmath__203_0_I3301 (.CO(inst_cellmath__203__W0[27]), .S(inst_cellmath__203__W1[26]), .A(N9879), .B(N8918), .CI(N9688));
XNOR2X1 inst_cellmath__203_0_I3302 (.Y(N9459), .A(N9736), .B(N9660));
OR2XL inst_cellmath__203_0_I3303 (.Y(N9841), .A(N9736), .B(N9660));
ADDFX1 inst_cellmath__203_0_I3304 (.CO(N9623), .S(N9230), .A(N9077), .B(N9459), .CI(N9386));
ADDFX1 inst_cellmath__203_0_I3305 (.CO(N8667), .S(N9987), .A(N10027), .B(N9231), .CI(N8937));
ADDFX1 inst_cellmath__203_0_I3306 (.CO(N9391), .S(N9008), .A(N10164), .B(N9884), .CI(N8694));
ADDFX1 inst_cellmath__203_0_I3307 (.CO(N10137), .S(N9780), .A(N9230), .B(N9431), .CI(N9987));
ADDFX1 inst_cellmath__203_0_I3308 (.CO(N9165), .S(N8796), .A(N9203), .B(N10172), .CI(N9008));
ADDFX1 inst_cellmath__203_0_I3309 (.CO(N9928), .S(N9557), .A(N9964), .B(N9780), .CI(N8796));
ADDFX1 inst_cellmath__203_0_I3310 (.CO(N8949), .S(N8613), .A(N9557), .B(N8981), .CI(N9751));
ADDFX1 inst_cellmath__203_0_I3311 (.CO(N9715), .S(N9329), .A(N8613), .B(N8769), .CI(N8770));
ADDFX1 inst_cellmath__203_0_I3312 (.CO(N8740), .S(N10073), .A(N8906), .B(N9083), .CI(N9274));
ADDFX1 inst_cellmath__203_0_I3313 (.CO(N9491), .S(N9098), .A(N9329), .B(N9466), .CI(N9525));
ADDFX1 inst_cellmath__203_0_I3314 (.CO(N10223), .S(N9869), .A(N10073), .B(N8592), .CI(N9098));
ADDFX1 inst_cellmath__203_0_I3315 (.CO(inst_cellmath__203__W0[28]), .S(inst_cellmath__203__W1[27]), .A(N10049), .B(N9296), .CI(N9869));
ADDFX1 inst_cellmath__203_0_I3317 (.CO(N10018), .S(N9654), .A(N9841), .B(N9315), .CI(N7288));
ADDFX1 inst_cellmath__203_0_I3318 (.CO(N9805), .S(N9425), .A(N8692), .B(N9621), .CI(N10237));
ADDFX1 inst_cellmath__203_0_I3319 (.CO(N8825), .S(N10163), .A(N9470), .B(N9772), .CI(N8826));
ADDFX1 inst_cellmath__203_0_I3320 (.CO(N9587), .S(N9194), .A(N9623), .B(N9654), .CI(N8667));
ADDFX1 inst_cellmath__203_0_I3321 (.CO(N8640), .S(N9955), .A(N9391), .B(N9425), .CI(N10163));
ADDFX1 inst_cellmath__203_0_I3322 (.CO(N9357), .S(N8973), .A(N10137), .B(N9194), .CI(N9955));
ADDFX1 inst_cellmath__203_0_I3323 (.CO(N10099), .S(N9744), .A(N8973), .B(N9165), .CI(N9928));
ADDFX1 inst_cellmath__203_0_I3324 (.CO(N9129), .S(N8765), .A(N8949), .B(N9744), .CI(N9404));
ADDFX1 inst_cellmath__203_0_I3325 (.CO(N9896), .S(N9519), .A(N8765), .B(N9523), .CI(N9475));
ADDFX1 inst_cellmath__203_0_I3326 (.CO(N8911), .S(N8587), .A(N9715), .B(N9666), .CI(N9849));
ADDFX1 inst_cellmath__203_0_I3327 (.CO(N9681), .S(N9289), .A(N9519), .B(N8740), .CI(N9491));
ADDFX1 inst_cellmath__203_0_I3328 (.CO(inst_cellmath__203__W0[29]), .S(inst_cellmath__203__W1[28]), .A(N10223), .B(N8587), .CI(N9289));
ADDFX1 inst_cellmath__203_0_I3329 (.CO(N9455), .S(N9063), .A(N9702), .B(N7390), .CI(N9040));
ADDFX1 inst_cellmath__203_0_I3330 (.CO(N10192), .S(N9832), .A(N9988), .B(N9195), .CI(N8901));
ADDFX1 inst_cellmath__203_0_I3331 (.CO(N9223), .S(N8849), .A(N10128), .B(N9851), .CI(N10018));
ADDFX1 inst_cellmath__203_0_I3332 (.CO(N9979), .S(N9615), .A(N8825), .B(N9805), .CI(N9063));
ADDFX1 inst_cellmath__203_0_I3333 (.CO(N9002), .S(N8661), .A(N9587), .B(N9832), .CI(N8849));
ADDFX1 inst_cellmath__203_0_I3334 (.CO(N9771), .S(N9385), .A(N8640), .B(N9615), .CI(N8661));
ADDFX1 inst_cellmath__203_0_I3335 (.CO(N8788), .S(N10130), .A(N9385), .B(N9357), .CI(N10099));
ADDFX1 inst_cellmath__203_0_I3336 (.CO(N9548), .S(N9157), .A(N8590), .B(N10130), .CI(N9129));
ADDFX1 inst_cellmath__203_0_I3337 (.CO(N8608), .S(N9919), .A(N10031), .B(N9856), .CI(N10203));
ADDFX1 inst_cellmath__203_0_I3338 (.CO(N9320), .S(N8942), .A(N9896), .B(N9157), .CI(N8911));
ADDFX1 inst_cellmath__203_0_I3339 (.CO(inst_cellmath__203__W0[30]), .S(inst_cellmath__203__W1[29]), .A(N9681), .B(N9919), .CI(N8942));
INVXL inst_cellmath__203_0_I3340 (.Y(N9362), .A(N9626));
ADDFX1 inst_cellmath__203_0_I3341 (.CO(N9091), .S(N8731), .A(N9588), .B(N9276), .CI(N9362));
ADDFX1 inst_cellmath__203_0_I3342 (.CO(N8875), .S(N10216), .A(N10206), .B(N8668), .CI(N9432));
ADDFX1 inst_cellmath__203_0_I3343 (.CO(N9644), .S(N9255), .A(N9455), .B(N8789), .CI(N10192));
ADDFX1 inst_cellmath__203_0_I3344 (.CO(N8678), .S(N10008), .A(N8731), .B(N9223), .CI(N10216));
ADDFX1 inst_cellmath__203_0_I3345 (.CO(N9415), .S(N9027), .A(N9255), .B(N9979), .CI(N9002));
ADDFX1 inst_cellmath__203_0_I3346 (.CO(N10158), .S(N9797), .A(N9771), .B(N10008), .CI(N9027));
ADDFX1 inst_cellmath__203_0_I3347 (.CO(N9186), .S(N8817), .A(N8788), .B(N9797), .CI(N9567));
ADDFX1 inst_cellmath__203_0_I3348 (.CO(N9946), .S(N9578), .A(N8817), .B(N9292), .CI(N8698));
ADDFX1 inst_cellmath__203_0_I3349 (.CO(N8967), .S(N8629), .A(N8863), .B(N9548), .CI(N8608));
ADDFX1 inst_cellmath__203_0_I3350 (.CO(inst_cellmath__203__W0[31]), .S(inst_cellmath__203__W1[30]), .A(N9320), .B(N9578), .CI(N8629));
ADDFX1 inst_cellmath__203_0_I3351 (.CO(N8758), .S(N10094), .A(N9668), .B(N9626), .CI(N9005));
ADDFX1 inst_cellmath__203_0_I3352 (.CO(N9510), .S(N9119), .A(N9956), .B(N9158), .CI(N8866));
ADDFX1 inst_cellmath__203_0_I3353 (.CO(N8579), .S(N9889), .A(N9091), .B(N9813), .CI(N8875));
ADDFX1 inst_cellmath__203_0_I3354 (.CO(N9283), .S(N8907), .A(N9119), .B(N10094), .CI(N9644));
ADDFX1 inst_cellmath__203_0_I3355 (.CO(N10038), .S(N9674), .A(N9889), .B(N8678), .CI(N8907));
ADDFX1 inst_cellmath__203_0_I3356 (.CO(N9056), .S(N8706), .A(N9674), .B(N9415), .CI(N10158));
ADDFX1 inst_cellmath__203_0_I3357 (.CO(N9824), .S(N9447), .A(N10047), .B(N8706), .CI(N9186));
ADDFX1 inst_cellmath__203_0_I3358 (.CO(N8845), .S(N10185), .A(N9238), .B(N9047), .CI(N9447));
ADDFX1 inst_cellmath__203_0_I3359 (.CO(inst_cellmath__203__W1[32]), .S(inst_cellmath__203__W1[31]), .A(N10185), .B(N9946), .CI(N8967));
INVXL inst_cellmath__203_0_I3360 (.Y(N9294), .A(N9785));
ADDFX1 inst_cellmath__203_0_I3361 (.CO(N8656), .S(N9974), .A(N9546), .B(N9242), .CI(N9294));
ADDFX1 inst_cellmath__203_0_I3362 (.CO(N10123), .S(N9763), .A(N10173), .B(N8638), .CI(N9392));
ADDFX1 inst_cellmath__203_0_I3363 (.CO(N9149), .S(N8782), .A(N9510), .B(N8758), .CI(N9974));
ADDFX1 inst_cellmath__203_0_I3364 (.CO(N9912), .S(N9539), .A(N8579), .B(N9763), .CI(N9283));
ADDFX1 inst_cellmath__203_0_I3365 (.CO(N8934), .S(N8601), .A(N9539), .B(N8782), .CI(N10038));
ADDFX1 inst_cellmath__203_0_I3366 (.CO(N9699), .S(N9311), .A(N9056), .B(N8601), .CI(N9066));
ADDFX1 inst_cellmath__203_0_I3367 (.CO(N8726), .S(N10061), .A(N9824), .B(N9723), .CI(N9311));
ADDFX1 inst_cellmath__203_0_I3368 (.CO(inst_cellmath__203__W1[33]), .S(inst_cellmath__203__W0[32]), .A(N10061), .B(N9627), .CI(N8845));
ADDFX1 inst_cellmath__203_0_I3369 (.CO(N10210), .S(N9854), .A(N9630), .B(N9785), .CI(N8974));
ADDFX1 inst_cellmath__203_0_I3370 (.CO(N9247), .S(N8870), .A(N8834), .B(N9920), .CI(N9781));
ADDFX1 inst_cellmath__203_0_I3371 (.CO(N10002), .S(N9637), .A(N10123), .B(N8656), .CI(N9854));
ADDFX1 inst_cellmath__203_0_I3372 (.CO(N9019), .S(N8674), .A(N9149), .B(N8870), .CI(N9637));
ADDFX1 inst_cellmath__203_0_I3373 (.CO(N9790), .S(N9407), .A(N8674), .B(N9912), .CI(N8934));
ADDFX1 inst_cellmath__203_0_I3374 (.CO(N8810), .S(N10150), .A(N9837), .B(N9407), .CI(N9699));
ADDFX1 inst_cellmath__203_0_I3375 (.CO(inst_cellmath__203__W1[34]), .S(inst_cellmath__203__W0[33]), .A(N10150), .B(N9996), .CI(N8726));
INVXL inst_cellmath__203_0_I3376 (.Y(N9228), .A(N9932));
ADDFX1 inst_cellmath__203_0_I3377 (.CO(N8624), .S(N9940), .A(N8609), .B(N9200), .CI(N9228));
ADDFX1 inst_cellmath__203_0_I3378 (.CO(N10088), .S(N9724), .A(N9358), .B(N10135), .CI(N10210));
ADDFX1 inst_cellmath__203_0_I3379 (.CO(N9109), .S(N8751), .A(N9940), .B(N9247), .CI(N9724));
ADDFX1 inst_cellmath__203_0_I3380 (.CO(N9883), .S(N9502), .A(N9019), .B(N10002), .CI(N8751));
ADDFX1 inst_cellmath__203_0_I3381 (.CO(N8897), .S(N10233), .A(N9790), .B(N9502), .CI(N8855));
ADDFX1 inst_cellmath__203_0_I3382 (.CO(inst_cellmath__203__W1[35]), .S(inst_cellmath__203__W0[34]), .A(N10233), .B(N9881), .CI(N8810));
ADDFX1 inst_cellmath__203_0_I3383 (.CO(N8699), .S(N10032), .A(N9595), .B(N9932), .CI(N8940));
ADDFX1 inst_cellmath__203_0_I3384 (.CO(N9438), .S(N9045), .A(N9742), .B(N8797), .CI(N8624));
ADDFX1 inst_cellmath__203_0_I3385 (.CO(N10178), .S(N9818), .A(N10088), .B(N10032), .CI(N9045));
ADDFX1 inst_cellmath__203_0_I3386 (.CO(N9208), .S(N8839), .A(N9818), .B(N9109), .CI(N9883));
ADDFX1 inst_cellmath__203_0_I3387 (.CO(inst_cellmath__203__W1[36]), .S(inst_cellmath__203__W0[35]), .A(N9620), .B(N8839), .CI(N8897));
INVXL inst_cellmath__203_0_I3388 (.Y(N9163), .A(N10077));
ADDFX1 inst_cellmath__203_0_I3389 (.CO(N8986), .S(N8648), .A(N10100), .B(N9166), .CI(N9163));
ADDFX1 inst_cellmath__203_0_I3390 (.CO(N8774), .S(N10114), .A(N8699), .B(N9321), .CI(N8648));
ADDFX1 inst_cellmath__203_0_I3391 (.CO(N9529), .S(N9140), .A(N10114), .B(N9438), .CI(N10178));
ADDFX1 inst_cellmath__203_0_I3392 (.CO(inst_cellmath__203__W1[37]), .S(inst_cellmath__203__W0[36]), .A(N9208), .B(N9140), .CI(N10121));
ADDFX1 inst_cellmath__203_0_I3393 (.CO(N9302), .S(N8924), .A(N9555), .B(N10077), .CI(N8766));
ADDFX1 inst_cellmath__203_0_I3394 (.CO(N10055), .S(N9691), .A(N8986), .B(N9707), .CI(N8924));
ADDFX1 inst_cellmath__203_0_I3395 (.CO(inst_cellmath__203__W1[38]), .S(inst_cellmath__203__W0[37]), .A(N9691), .B(N8774), .CI(N9529));
ADDFX1 inst_cellmath__203_0_I3396 (.CO(N9847), .S(N9467), .A(N9128), .B(N10228), .CI(N10066));
ADDFX1 inst_cellmath__203_0_I3397 (.CO(inst_cellmath__203__W1[39]), .S(inst_cellmath__203__W0[38]), .A(N9467), .B(N9302), .CI(N10055));
INVXL inst_cellmath__203_0_I3398 (.Y(N9236), .A(N9628));
ADDFX1 inst_cellmath__203_0_I3399 (.CO(inst_cellmath__203__W1[40]), .S(inst_cellmath__203__W0[39]), .A(N8732), .B(N9236), .CI(N9847));
ADDFX1 inst_cellmath__203_0_I3400 (.CO(inst_cellmath__203__W1[41]), .S(inst_cellmath__203__W0[40]), .A(N9628), .B(N8689), .CI(N9092));
INVXL inst_cellmath__203_0_I3401 (.Y(inst_cellmath__203__W0[41]), .A(inst_cellmath__203__W1[42]));
ADDHX1 cynw_cm_float_cos_I3404 (.CO(N12044), .S(N11910), .A(inst_cellmath__195[0]), .B(inst_cellmath__203__W0[18]));
ADDFX1 cynw_cm_float_cos_I3405 (.CO(N12322), .S(N12183), .A(inst_cellmath__203__W0[19]), .B(inst_cellmath__195[1]), .CI(inst_cellmath__203__W1[19]));
ADDFX1 cynw_cm_float_cos_I3406 (.CO(N11965), .S(N11833), .A(inst_cellmath__203__W0[20]), .B(inst_cellmath__195[2]), .CI(inst_cellmath__203__W1[20]));
ADDFX1 cynw_cm_float_cos_I3407 (.CO(N12238), .S(N12104), .A(inst_cellmath__203__W0[21]), .B(inst_cellmath__195[3]), .CI(inst_cellmath__203__W1[21]));
ADDFX1 cynw_cm_float_cos_I3408 (.CO(N11886), .S(N12382), .A(inst_cellmath__203__W0[22]), .B(inst_cellmath__195[4]), .CI(inst_cellmath__203__W1[22]));
ADDFX1 cynw_cm_float_cos_I3409 (.CO(N12160), .S(N12019), .A(inst_cellmath__203__W0[23]), .B(inst_cellmath__195[5]), .CI(inst_cellmath__203__W1[23]));
ADDFX1 cynw_cm_float_cos_I3410 (.CO(N12435), .S(N12299), .A(inst_cellmath__203__W0[24]), .B(inst_cellmath__195[6]), .CI(inst_cellmath__203__W1[24]));
ADDFX1 cynw_cm_float_cos_I3411 (.CO(N12079), .S(N11943), .A(inst_cellmath__203__W0[25]), .B(inst_cellmath__195[7]), .CI(inst_cellmath__203__W1[25]));
ADDFX1 cynw_cm_float_cos_I3412 (.CO(N12358), .S(N12215), .A(inst_cellmath__203__W0[26]), .B(inst_cellmath__195[8]), .CI(inst_cellmath__203__W1[26]));
ADDFX1 cynw_cm_float_cos_I3413 (.CO(N11995), .S(N11864), .A(inst_cellmath__203__W0[27]), .B(inst_cellmath__195[9]), .CI(inst_cellmath__203__W1[27]));
ADDFX1 cynw_cm_float_cos_I3414 (.CO(N12276), .S(N12137), .A(inst_cellmath__203__W0[28]), .B(inst_cellmath__195[10]), .CI(inst_cellmath__203__W1[28]));
ADDFX1 cynw_cm_float_cos_I3415 (.CO(N11921), .S(N12413), .A(inst_cellmath__203__W0[29]), .B(inst_cellmath__195[11]), .CI(inst_cellmath__203__W1[29]));
ADDFX1 cynw_cm_float_cos_I3416 (.CO(N12193), .S(N12055), .A(inst_cellmath__203__W0[30]), .B(inst_cellmath__195[12]), .CI(inst_cellmath__203__W1[30]));
ADDFX1 cynw_cm_float_cos_I3417 (.CO(N11844), .S(N12335), .A(inst_cellmath__203__W0[31]), .B(inst_cellmath__195[13]), .CI(inst_cellmath__203__W1[31]));
ADDFX1 cynw_cm_float_cos_I3418 (.CO(N12116), .S(N11976), .A(inst_cellmath__203__W0[32]), .B(inst_cellmath__195[14]), .CI(inst_cellmath__203__W1[32]));
ADDFX1 cynw_cm_float_cos_I3419 (.CO(N12393), .S(N12251), .A(inst_cellmath__203__W1[33]), .B(inst_cellmath__195[15]), .CI(inst_cellmath__203__W0[33]));
ADDFX1 cynw_cm_float_cos_I3420 (.CO(N12032), .S(N11897), .A(inst_cellmath__203__W0[34]), .B(inst_cellmath__195[16]), .CI(inst_cellmath__203__W1[34]));
ADDFX1 cynw_cm_float_cos_I3421 (.CO(N12311), .S(N12171), .A(inst_cellmath__203__W1[35]), .B(inst_cellmath__195[17]), .CI(inst_cellmath__203__W0[35]));
ADDFX1 cynw_cm_float_cos_I3422 (.CO(N11953), .S(N12449), .A(inst_cellmath__203__W0[36]), .B(inst_cellmath__195[18]), .CI(inst_cellmath__203__W1[36]));
ADDFX1 cynw_cm_float_cos_I3423 (.CO(N12225), .S(N12091), .A(inst_cellmath__203__W0[37]), .B(inst_cellmath__195[19]), .CI(inst_cellmath__203__W1[37]));
ADDFX1 cynw_cm_float_cos_I3424 (.CO(N11873), .S(N12370), .A(inst_cellmath__203__W0[38]), .B(inst_cellmath__195[20]), .CI(inst_cellmath__203__W1[38]));
ADDFX1 cynw_cm_float_cos_I3425 (.CO(N12147), .S(N12007), .A(inst_cellmath__203__W0[39]), .B(inst_cellmath__195[21]), .CI(inst_cellmath__203__W1[39]));
ADDFX1 cynw_cm_float_cos_I3426 (.CO(N12422), .S(N12287), .A(inst_cellmath__203__W0[40]), .B(inst_cellmath__195[22]), .CI(inst_cellmath__203__W1[40]));
ADDFX1 cynw_cm_float_cos_I3427 (.CO(N12066), .S(N11931), .A(inst_cellmath__195[23]), .B(inst_cellmath__203__W0[41]), .CI(inst_cellmath__203__W1[41]));
ADDFX1 cynw_cm_float_cos_I3428 (.CO(N12344), .S(N12204), .A(inst_cellmath__203__W1[42]), .B(inst_cellmath__203__W0[42]), .CI(inst_cellmath__195[24]));
ADDHX1 cynw_cm_float_cos_I3429 (.CO(N11983), .S(N11853), .A(1'B1), .B(inst_cellmath__195[25]));
ADDHX1 cynw_cm_float_cos_I3430 (.CO(N12262), .S(N12122), .A(1'B1), .B(inst_cellmath__195[26]));
ADDHX1 cynw_cm_float_cos_I3431 (.CO(N11904), .S(N12399), .A(1'B1), .B(inst_cellmath__195[27]));
INVXL hap1_A_I23530 (.Y(N12042), .A(inst_cellmath__195[28]));
OR2XL hap1_A_I8389 (.Y(N12178), .A(1'B0), .B(inst_cellmath__195[28]));
AND2XL cynw_cm_float_cos_I8339 (.Y(N12317), .A(N6554), .B(N6280));
AND2XL cynw_cm_float_cos_I3438 (.Y(N12155), .A(inst_cellmath__203__W0[2]), .B(inst_cellmath__203__W1[2]));
NOR2XL cynw_cm_float_cos_I3439 (.Y(N12295), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
NAND2XL cynw_cm_float_cos_I3440 (.Y(N12433), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
AND2XL cynw_cm_float_cos_I3442 (.Y(N12075), .A(inst_cellmath__203__W0[4]), .B(inst_cellmath__203__W1[4]));
NOR2XL cynw_cm_float_cos_I3443 (.Y(N12213), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
NAND2XL cynw_cm_float_cos_I3444 (.Y(N12353), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
AND2XL cynw_cm_float_cos_I3446 (.Y(N11993), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
NOR2XL cynw_cm_float_cos_I3447 (.Y(N12130), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
NAND2XL cynw_cm_float_cos_I3448 (.Y(N12272), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
AND2XL cynw_cm_float_cos_I3450 (.Y(N11916), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
NOR2XL cynw_cm_float_cos_I3451 (.Y(N12051), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
NAND2XL cynw_cm_float_cos_I3452 (.Y(N12191), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
AND2XL cynw_cm_float_cos_I3454 (.Y(N11840), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
NOR2XL cynw_cm_float_cos_I3455 (.Y(N11974), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
NAND2XL cynw_cm_float_cos_I3456 (.Y(N12112), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
AND2XL cynw_cm_float_cos_I3458 (.Y(N12391), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
NOR2XL cynw_cm_float_cos_I3459 (.Y(N11893), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NAND2XL cynw_cm_float_cos_I3460 (.Y(N12028), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NOR2XL cynw_cm_float_cos_I3461 (.Y(N12169), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NAND2XL cynw_cm_float_cos_I3462 (.Y(N12307), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NOR2XL cynw_cm_float_cos_I3463 (.Y(N12445), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NOR2XL cynw_cm_float_cos_I3465 (.Y(N12087), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
NAND2XL cynw_cm_float_cos_I3466 (.Y(N12223), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
NOR2XL cynw_cm_float_cos_I3467 (.Y(N12368), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NOR2XL cynw_cm_float_cos_I3469 (.Y(N12005), .A(inst_cellmath__203__W1[18]), .B(N11910));
NAND2XL cynw_cm_float_cos_I3470 (.Y(N12145), .A(inst_cellmath__203__W1[18]), .B(N11910));
NOR2XL cynw_cm_float_cos_I3471 (.Y(N12283), .A(N12044), .B(N12183));
NAND2XL cynw_cm_float_cos_I3472 (.Y(N12419), .A(N12044), .B(N12183));
AND2XL cynw_cm_float_cos_I23531 (.Y(N12201), .A(inst_cellmath__203__W0[1]), .B(inst_cellmath__203__W1[1]));
OAI22XL cynw_cm_float_cos_I8340 (.Y(N12037), .A0(N12155), .A1(N12201), .B0(inst_cellmath__203__W0[2]), .B1(inst_cellmath__203__W1[2]));
AOI21XL cynw_cm_float_cos_I3477 (.Y(N11879), .A0(N12433), .A1(N12037), .B0(N12295));
OAI22XL cynw_cm_float_cos_I8341 (.Y(N12269), .A0(N12075), .A1(N11879), .B0(inst_cellmath__203__W0[4]), .B1(inst_cellmath__203__W1[4]));
AOI21XL cynw_cm_float_cos_I3481 (.Y(N12025), .A0(N12353), .A1(N12269), .B0(N12213));
OAI22XL cynw_cm_float_cos_I8342 (.Y(N12340), .A0(N11993), .A1(N12025), .B0(inst_cellmath__203__W0[6]), .B1(inst_cellmath__203__W1[6]));
AOI21XL cynw_cm_float_cos_I3485 (.Y(N12011), .A0(N12272), .A1(N12340), .B0(N12130));
OAI22XL cynw_cm_float_cos_I8343 (.Y(N12241), .A0(N11916), .A1(N12011), .B0(inst_cellmath__203__W0[8]), .B1(inst_cellmath__203__W1[8]));
AOI21XL cynw_cm_float_cos_I3489 (.Y(N11847), .A0(N12191), .A1(N12241), .B0(N12051));
OAI22XL cynw_cm_float_cos_I8344 (.Y(N11986), .A0(N11840), .A1(N11847), .B0(inst_cellmath__203__W0[10]), .B1(inst_cellmath__203__W1[10]));
AOI21XL cynw_cm_float_cos_I3493 (.Y(N12134), .A0(N12112), .A1(N11986), .B0(N11974));
OAI22XL cynw_cm_float_cos_I8345 (.Y(N12203), .A0(N12391), .A1(N12134), .B0(inst_cellmath__203__W0[12]), .B1(inst_cellmath__203__W1[12]));
AO21XL cynw_cm_float_cos_I3497 (.Y(N12425), .A0(N12307), .A1(N11893), .B0(N12169));
AOI31X1 cynw_cm_float_cos_I3499 (.Y(N12388), .A0(N12307), .A1(N12028), .A2(N12203), .B0(N12425));
AOI21XL cynw_cm_float_cos_I3500 (.Y(N12305), .A0(N12223), .A1(N12445), .B0(N12087));
OAI2BB1X1 cynw_cm_float_cos_I8346 (.Y(N12443), .A0N(inst_cellmath__203__W0[15]), .A1N(inst_cellmath__203__W1[15]), .B0(N12223));
AOI21XL cynw_cm_float_cos_I3503 (.Y(N12221), .A0(N12145), .A1(N12368), .B0(N12005));
OAI2BB1X1 cynw_cm_float_cos_I8347 (.Y(N12365), .A0N(inst_cellmath__203__W0[17]), .A1N(inst_cellmath__203__W1[17]), .B0(N12145));
OAI21XL cynw_cm_float_cos_I3508 (.Y(N11900), .A0(N12365), .A1(N12305), .B0(N12221));
NOR3XL cynw_cm_float_cos_I3509 (.Y(N12254), .A(N12365), .B(N12443), .C(N12388));
OR2XL cynw_cm_float_cos_I3510 (.Y(N12082), .A(N12254), .B(N11900));
AO21XL cynw_cm_float_cos_I3554 (.Y(N12062), .A0(N12419), .A1(N12082), .B0(N12283));
NOR2XL cynw_cm_float_cos_I3555 (.Y(N12343), .A(N12322), .B(N11833));
NAND2XL cynw_cm_float_cos_I3556 (.Y(N11850), .A(N12322), .B(N11833));
NOR2XL cynw_cm_float_cos_I3557 (.Y(N11980), .A(N11965), .B(N12104));
NAND2XL cynw_cm_float_cos_I3558 (.Y(N12121), .A(N11965), .B(N12104));
NOR2XL cynw_cm_float_cos_I3559 (.Y(N12257), .A(N12238), .B(N12382));
NAND2XL cynw_cm_float_cos_I3560 (.Y(N12396), .A(N12238), .B(N12382));
NOR2XL cynw_cm_float_cos_I3561 (.Y(N11903), .A(N11886), .B(N12019));
NAND2XL cynw_cm_float_cos_I3562 (.Y(N12038), .A(N11886), .B(N12019));
NOR2XL cynw_cm_float_cos_I3563 (.Y(N12175), .A(N12160), .B(N12299));
NAND2XL cynw_cm_float_cos_I3564 (.Y(N12316), .A(N12160), .B(N12299));
NOR2XL cynw_cm_float_cos_I3565 (.Y(N11827), .A(N12435), .B(N11943));
NAND2XL cynw_cm_float_cos_I3566 (.Y(N11958), .A(N12435), .B(N11943));
NOR2XL cynw_cm_float_cos_I3567 (.Y(N12099), .A(N12079), .B(N12215));
NAND2XL cynw_cm_float_cos_I3568 (.Y(N12232), .A(N12079), .B(N12215));
NOR2XL cynw_cm_float_cos_I3569 (.Y(N12374), .A(N12358), .B(N11864));
NAND2XL cynw_cm_float_cos_I3570 (.Y(N11880), .A(N12358), .B(N11864));
NOR2XL cynw_cm_float_cos_I3571 (.Y(N12014), .A(N11995), .B(N12137));
NAND2XL cynw_cm_float_cos_I3572 (.Y(N12152), .A(N11995), .B(N12137));
NOR2XL cynw_cm_float_cos_I3573 (.Y(N12293), .A(N12276), .B(N12413));
NAND2XL cynw_cm_float_cos_I3574 (.Y(N12430), .A(N12276), .B(N12413));
NOR2XL cynw_cm_float_cos_I3575 (.Y(N11935), .A(N11921), .B(N12055));
NAND2XL cynw_cm_float_cos_I3576 (.Y(N12073), .A(N11921), .B(N12055));
NOR2XL cynw_cm_float_cos_I3577 (.Y(N12210), .A(N12193), .B(N12335));
NAND2XL cynw_cm_float_cos_I3578 (.Y(N12350), .A(N12193), .B(N12335));
NOR2XL cynw_cm_float_cos_I3579 (.Y(N11858), .A(N11844), .B(N11976));
NAND2XL cynw_cm_float_cos_I3580 (.Y(N11990), .A(N11844), .B(N11976));
NOR2XL cynw_cm_float_cos_I3581 (.Y(N12127), .A(N12116), .B(N12251));
NAND2XL cynw_cm_float_cos_I3582 (.Y(N12270), .A(N12116), .B(N12251));
NOR2XL cynw_cm_float_cos_I3583 (.Y(N12408), .A(N12393), .B(N11897));
NAND2XL cynw_cm_float_cos_I3584 (.Y(N11913), .A(N12393), .B(N11897));
NOR2XL cynw_cm_float_cos_I3585 (.Y(N12049), .A(N12032), .B(N12171));
NAND2XL cynw_cm_float_cos_I3586 (.Y(N12188), .A(N12032), .B(N12171));
NOR2XL cynw_cm_float_cos_I3587 (.Y(N12327), .A(N12449), .B(N12311));
NAND2XL cynw_cm_float_cos_I3588 (.Y(N11838), .A(N12449), .B(N12311));
NOR2XL cynw_cm_float_cos_I3589 (.Y(N11971), .A(N12091), .B(N11953));
NAND2XL cynw_cm_float_cos_I3590 (.Y(N12108), .A(N12091), .B(N11953));
NOR2XL cynw_cm_float_cos_I3591 (.Y(N12245), .A(N12370), .B(N12225));
NAND2XL cynw_cm_float_cos_I3592 (.Y(N12387), .A(N12370), .B(N12225));
NOR2XL cynw_cm_float_cos_I3593 (.Y(N11890), .A(N12007), .B(N11873));
NAND2XL cynw_cm_float_cos_I3594 (.Y(N12026), .A(N12007), .B(N11873));
NOR2XL cynw_cm_float_cos_I3595 (.Y(N12166), .A(N12287), .B(N12147));
NAND2XL cynw_cm_float_cos_I3596 (.Y(N12303), .A(N12287), .B(N12147));
NOR2XL cynw_cm_float_cos_I3597 (.Y(N12442), .A(N11931), .B(N12422));
NAND2XL cynw_cm_float_cos_I3598 (.Y(N11948), .A(N11931), .B(N12422));
NOR2XL cynw_cm_float_cos_I3599 (.Y(N12084), .A(N12204), .B(N12066));
NAND2XL cynw_cm_float_cos_I3600 (.Y(N12220), .A(N12204), .B(N12066));
NOR2XL cynw_cm_float_cos_I3601 (.Y(N12364), .A(N12344), .B(N11853));
NAND2XL cynw_cm_float_cos_I3602 (.Y(N11867), .A(N12344), .B(N11853));
NOR2XL cynw_cm_float_cos_I3603 (.Y(N12002), .A(N11983), .B(N12122));
NAND2XL cynw_cm_float_cos_I3604 (.Y(N12142), .A(N11983), .B(N12122));
NOR2XL cynw_cm_float_cos_I3605 (.Y(N12281), .A(N12262), .B(N12399));
NAND2XL cynw_cm_float_cos_I3606 (.Y(N12418), .A(N12262), .B(N12399));
NOR2XL cynw_cm_float_cos_I3607 (.Y(N11928), .A(N12042), .B(N11904));
NAND2XL cynw_cm_float_cos_I3608 (.Y(N12059), .A(N12042), .B(N11904));
NOR2XL cynw_cm_float_cos_I3609 (.Y(N12200), .A(N12317), .B(N12178));
NAND2XL cynw_cm_float_cos_I3610 (.Y(N12341), .A(N12317), .B(N12178));
AO21XL cynw_cm_float_cos_I3611 (.Y(N12255), .A0(N11850), .A1(N12062), .B0(N12343));
AO21XL cynw_cm_float_cos_I3612 (.Y(N11901), .A0(N12121), .A1(N12343), .B0(N11980));
AND2XL cynw_cm_float_cos_I3613 (.Y(N12035), .A(N12121), .B(N11850));
AO21XL cynw_cm_float_cos_I3614 (.Y(N12174), .A0(N12396), .A1(N11980), .B0(N12257));
AND2XL cynw_cm_float_cos_I3615 (.Y(N12314), .A(N12396), .B(N12121));
AO21XL cynw_cm_float_cos_I3616 (.Y(N12452), .A0(N12038), .A1(N12257), .B0(N11903));
AND2XL cynw_cm_float_cos_I3617 (.Y(N11956), .A(N12038), .B(N12396));
AO21XL cynw_cm_float_cos_I3618 (.Y(N12097), .A0(N12316), .A1(N11903), .B0(N12175));
AND2XL cynw_cm_float_cos_I3619 (.Y(N12228), .A(N12316), .B(N12038));
AO21XL cynw_cm_float_cos_I3620 (.Y(N12373), .A0(N11958), .A1(N12175), .B0(N11827));
AND2XL cynw_cm_float_cos_I3621 (.Y(N11876), .A(N11958), .B(N12316));
AO21XL cynw_cm_float_cos_I3622 (.Y(N12012), .A0(N12232), .A1(N11827), .B0(N12099));
AND2XL cynw_cm_float_cos_I3623 (.Y(N12150), .A(N12232), .B(N11958));
AO21XL cynw_cm_float_cos_I3624 (.Y(N12291), .A0(N11880), .A1(N12099), .B0(N12374));
AND2XL cynw_cm_float_cos_I3625 (.Y(N12427), .A(N11880), .B(N12232));
AO21XL cynw_cm_float_cos_I3626 (.Y(N11934), .A0(N12152), .A1(N12374), .B0(N12014));
AND2XL cynw_cm_float_cos_I3627 (.Y(N12070), .A(N12152), .B(N11880));
AO21XL cynw_cm_float_cos_I3628 (.Y(N12208), .A0(N12430), .A1(N12014), .B0(N12293));
AND2XL cynw_cm_float_cos_I3629 (.Y(N12348), .A(N12430), .B(N12152));
AO21XL cynw_cm_float_cos_I3630 (.Y(N11856), .A0(N12073), .A1(N12293), .B0(N11935));
AND2XL cynw_cm_float_cos_I3631 (.Y(N11988), .A(N12073), .B(N12430));
AO21XL cynw_cm_float_cos_I3632 (.Y(N12126), .A0(N12350), .A1(N11935), .B0(N12210));
AND2XL cynw_cm_float_cos_I3633 (.Y(N12267), .A(N12350), .B(N12073));
AO21XL cynw_cm_float_cos_I3634 (.Y(N12405), .A0(N11990), .A1(N12210), .B0(N11858));
AND2XL cynw_cm_float_cos_I3635 (.Y(N11911), .A(N11990), .B(N12350));
AO21XL cynw_cm_float_cos_I3636 (.Y(N12047), .A0(N12270), .A1(N11858), .B0(N12127));
AND2XL cynw_cm_float_cos_I3637 (.Y(N12184), .A(N12270), .B(N11990));
AO21XL cynw_cm_float_cos_I3638 (.Y(N12325), .A0(N11913), .A1(N12127), .B0(N12408));
AND2XL cynw_cm_float_cos_I3639 (.Y(N11836), .A(N11913), .B(N12270));
AO21XL cynw_cm_float_cos_I3640 (.Y(N11967), .A0(N12188), .A1(N12408), .B0(N12049));
AND2XL cynw_cm_float_cos_I3641 (.Y(N12105), .A(N12188), .B(N11913));
AO21XL cynw_cm_float_cos_I3642 (.Y(N12243), .A0(N11838), .A1(N12049), .B0(N12327));
AND2XL cynw_cm_float_cos_I3643 (.Y(N12383), .A(N11838), .B(N12188));
AO21XL cynw_cm_float_cos_I3644 (.Y(N11888), .A0(N12108), .A1(N12327), .B0(N11971));
AND2XL cynw_cm_float_cos_I3645 (.Y(N12023), .A(N12108), .B(N11838));
AO21XL cynw_cm_float_cos_I3646 (.Y(N12162), .A0(N12387), .A1(N11971), .B0(N12245));
AND2XL cynw_cm_float_cos_I3647 (.Y(N12300), .A(N12387), .B(N12108));
AO21XL cynw_cm_float_cos_I3648 (.Y(N12439), .A0(N12026), .A1(N12245), .B0(N11890));
AND2XL cynw_cm_float_cos_I3649 (.Y(N11944), .A(N12026), .B(N12387));
AO21XL cynw_cm_float_cos_I3650 (.Y(N12081), .A0(N12303), .A1(N11890), .B0(N12166));
AND2XL cynw_cm_float_cos_I3651 (.Y(N12218), .A(N12303), .B(N12026));
AO21XL cynw_cm_float_cos_I3652 (.Y(N12360), .A0(N11948), .A1(N12166), .B0(N12442));
AND2XL cynw_cm_float_cos_I3653 (.Y(N11865), .A(N11948), .B(N12303));
AO21XL cynw_cm_float_cos_I3654 (.Y(N12000), .A0(N12220), .A1(N12442), .B0(N12084));
AND2XL cynw_cm_float_cos_I3655 (.Y(N12138), .A(N12220), .B(N11948));
AO21XL cynw_cm_float_cos_I3656 (.Y(N12278), .A0(N11867), .A1(N12084), .B0(N12364));
AND2XL cynw_cm_float_cos_I3657 (.Y(N12416), .A(N11867), .B(N12220));
AO21XL cynw_cm_float_cos_I3658 (.Y(N11923), .A0(N12142), .A1(N12364), .B0(N12002));
AND2XL cynw_cm_float_cos_I3659 (.Y(N12056), .A(N12142), .B(N11867));
AO21XL cynw_cm_float_cos_I3660 (.Y(N12198), .A0(N12418), .A1(N12002), .B0(N12281));
AND2XL cynw_cm_float_cos_I3661 (.Y(N12336), .A(N12418), .B(N12142));
AO21XL cynw_cm_float_cos_I3662 (.Y(N11848), .A0(N12059), .A1(N12281), .B0(N11928));
AND2XL cynw_cm_float_cos_I3663 (.Y(N11979), .A(N12059), .B(N12418));
AO21XL cynw_cm_float_cos_I3664 (.Y(N12117), .A0(N12341), .A1(N11928), .B0(N12200));
AND2XL cynw_cm_float_cos_I3665 (.Y(N12253), .A(N12341), .B(N12059));
AND2XL cynw_cm_float_cos_I3666 (.Y(N12034), .A(N12317), .B(N12341));
AO21XL cynw_cm_float_cos_I3667 (.Y(N12092), .A0(N12035), .A1(N12062), .B0(N11901));
AO21XL cynw_cm_float_cos_I3668 (.Y(N12372), .A0(N12314), .A1(N12255), .B0(N12174));
AO21XL cynw_cm_float_cos_I3669 (.Y(N12010), .A0(N11956), .A1(N11901), .B0(N12452));
AND2XL cynw_cm_float_cos_I3670 (.Y(N12149), .A(N11956), .B(N12035));
AO21XL cynw_cm_float_cos_I3671 (.Y(N12288), .A0(N12228), .A1(N12174), .B0(N12097));
AND2XL cynw_cm_float_cos_I3672 (.Y(N12426), .A(N12228), .B(N12314));
AO21XL cynw_cm_float_cos_I3673 (.Y(N11933), .A0(N11876), .A1(N12452), .B0(N12373));
AND2XL cynw_cm_float_cos_I3674 (.Y(N12068), .A(N11876), .B(N11956));
AO21XL cynw_cm_float_cos_I3675 (.Y(N12207), .A0(N12150), .A1(N12097), .B0(N12012));
AND2XL cynw_cm_float_cos_I3676 (.Y(N12347), .A(N12150), .B(N12228));
AO21XL cynw_cm_float_cos_I3677 (.Y(N11854), .A0(N12427), .A1(N12373), .B0(N12291));
AND2XL cynw_cm_float_cos_I3678 (.Y(N11987), .A(N12427), .B(N11876));
AO21XL cynw_cm_float_cos_I3679 (.Y(N12125), .A0(N12070), .A1(N12012), .B0(N11934));
AND2XL cynw_cm_float_cos_I3680 (.Y(N12265), .A(N12070), .B(N12150));
AO21XL cynw_cm_float_cos_I3681 (.Y(N12403), .A0(N12348), .A1(N12291), .B0(N12208));
AND2XL cynw_cm_float_cos_I3682 (.Y(N11909), .A(N12348), .B(N12427));
AO21XL cynw_cm_float_cos_I3683 (.Y(N12045), .A0(N11988), .A1(N11934), .B0(N11856));
AND2XL cynw_cm_float_cos_I3684 (.Y(N12182), .A(N11988), .B(N12070));
AO21XL cynw_cm_float_cos_I3685 (.Y(N12321), .A0(N12267), .A1(N12208), .B0(N12126));
AND2XL cynw_cm_float_cos_I3686 (.Y(N11834), .A(N12267), .B(N12348));
AO21XL cynw_cm_float_cos_I3687 (.Y(N11964), .A0(N11911), .A1(N11856), .B0(N12405));
AND2XL cynw_cm_float_cos_I3688 (.Y(N12103), .A(N11911), .B(N11988));
AO21XL cynw_cm_float_cos_I3689 (.Y(N12239), .A0(N12184), .A1(N12126), .B0(N12047));
AND2XL cynw_cm_float_cos_I3690 (.Y(N12381), .A(N12184), .B(N12267));
AO21XL cynw_cm_float_cos_I3691 (.Y(N11885), .A0(N11836), .A1(N12405), .B0(N12325));
AND2XL cynw_cm_float_cos_I3692 (.Y(N12021), .A(N11836), .B(N11911));
AO21XL cynw_cm_float_cos_I3693 (.Y(N12159), .A0(N12105), .A1(N12047), .B0(N11967));
AND2XL cynw_cm_float_cos_I3694 (.Y(N12298), .A(N12105), .B(N12184));
AO21XL cynw_cm_float_cos_I3695 (.Y(N12436), .A0(N12383), .A1(N12325), .B0(N12243));
AND2XL cynw_cm_float_cos_I3696 (.Y(N11942), .A(N12383), .B(N11836));
AO21XL cynw_cm_float_cos_I3697 (.Y(N12078), .A0(N12023), .A1(N11967), .B0(N11888));
AND2XL cynw_cm_float_cos_I3698 (.Y(N12216), .A(N12023), .B(N12105));
AO21XL cynw_cm_float_cos_I3699 (.Y(N12357), .A0(N12300), .A1(N12243), .B0(N12162));
AND2XL cynw_cm_float_cos_I3700 (.Y(N11863), .A(N12300), .B(N12383));
AO21XL cynw_cm_float_cos_I3701 (.Y(N11997), .A0(N11944), .A1(N11888), .B0(N12439));
AND2XL cynw_cm_float_cos_I3702 (.Y(N12136), .A(N11944), .B(N12023));
AO21XL cynw_cm_float_cos_I3703 (.Y(N12275), .A0(N12218), .A1(N12162), .B0(N12081));
AND2XL cynw_cm_float_cos_I3704 (.Y(N12414), .A(N12218), .B(N12300));
AO21XL cynw_cm_float_cos_I3705 (.Y(N11920), .A0(N11865), .A1(N12439), .B0(N12360));
AND2XL cynw_cm_float_cos_I3706 (.Y(N12054), .A(N11865), .B(N11944));
AO21XL cynw_cm_float_cos_I3707 (.Y(N12194), .A0(N12138), .A1(N12081), .B0(N12000));
AND2XL cynw_cm_float_cos_I3708 (.Y(N12334), .A(N12138), .B(N12218));
AO21XL cynw_cm_float_cos_I3709 (.Y(N11843), .A0(N12416), .A1(N12360), .B0(N12278));
AND2XL cynw_cm_float_cos_I3710 (.Y(N11977), .A(N12416), .B(N11865));
AO21XL cynw_cm_float_cos_I3711 (.Y(N12115), .A0(N12056), .A1(N12000), .B0(N11923));
AND2XL cynw_cm_float_cos_I3712 (.Y(N12250), .A(N12056), .B(N12138));
AO21XL cynw_cm_float_cos_I3713 (.Y(N12394), .A0(N12336), .A1(N12278), .B0(N12198));
AND2XL cynw_cm_float_cos_I3714 (.Y(N11896), .A(N12336), .B(N12416));
AO21XL cynw_cm_float_cos_I3715 (.Y(N12031), .A0(N11979), .A1(N11923), .B0(N11848));
AND2XL cynw_cm_float_cos_I3716 (.Y(N12172), .A(N11979), .B(N12056));
AO21XL cynw_cm_float_cos_I3717 (.Y(N12310), .A0(N12253), .A1(N12198), .B0(N12117));
AND2XL cynw_cm_float_cos_I3718 (.Y(N12448), .A(N12253), .B(N12336));
AO22XL cynw_cm_float_cos_I3719 (.Y(N11954), .A0(N12317), .A1(N12200), .B0(N12034), .B1(N11848));
AND2XL cynw_cm_float_cos_I3720 (.Y(N12090), .A(N12034), .B(N11979));
AO21XL cynw_cm_float_cos_I3721 (.Y(N12065), .A0(N12149), .A1(N12062), .B0(N12010));
AO21XL cynw_cm_float_cos_I3722 (.Y(N12345), .A0(N12426), .A1(N12255), .B0(N12288));
AO21XL cynw_cm_float_cos_I3723 (.Y(N11982), .A0(N12068), .A1(N12092), .B0(N11933));
AO21XL cynw_cm_float_cos_I3724 (.Y(N12261), .A0(N12347), .A1(N12372), .B0(N12207));
AO21XL cynw_cm_float_cos_I3725 (.Y(N11906), .A0(N11987), .A1(N12010), .B0(N11854));
AND2XL cynw_cm_float_cos_I3726 (.Y(N12041), .A(N11987), .B(N12149));
AO21XL cynw_cm_float_cos_I3727 (.Y(N12177), .A0(N12265), .A1(N12288), .B0(N12125));
AND2XL cynw_cm_float_cos_I3728 (.Y(N12318), .A(N12265), .B(N12426));
AO21XL cynw_cm_float_cos_I3729 (.Y(N11830), .A0(N11909), .A1(N11933), .B0(N12403));
AND2XL cynw_cm_float_cos_I3730 (.Y(N11960), .A(N11909), .B(N12068));
AO21XL cynw_cm_float_cos_I3731 (.Y(N12100), .A0(N12182), .A1(N12207), .B0(N12045));
AND2XL cynw_cm_float_cos_I3732 (.Y(N12235), .A(N12182), .B(N12347));
AO21XL cynw_cm_float_cos_I3733 (.Y(N12376), .A0(N11834), .A1(N11854), .B0(N12321));
AND2XL cynw_cm_float_cos_I3734 (.Y(N11881), .A(N11834), .B(N11987));
AO21XL cynw_cm_float_cos_I3735 (.Y(N12016), .A0(N12103), .A1(N12125), .B0(N11964));
AND2XL cynw_cm_float_cos_I3736 (.Y(N12154), .A(N12103), .B(N12265));
AO21XL cynw_cm_float_cos_I3737 (.Y(N12294), .A0(N12381), .A1(N12403), .B0(N12239));
AND2XL cynw_cm_float_cos_I3738 (.Y(N12432), .A(N12381), .B(N11909));
AO21XL cynw_cm_float_cos_I3739 (.Y(N11937), .A0(N12021), .A1(N12045), .B0(N11885));
AND2XL cynw_cm_float_cos_I3740 (.Y(N12074), .A(N12021), .B(N12182));
AO21XL cynw_cm_float_cos_I3741 (.Y(N12212), .A0(N12298), .A1(N12321), .B0(N12159));
AND2XL cynw_cm_float_cos_I3742 (.Y(N12352), .A(N12298), .B(N11834));
AO21XL cynw_cm_float_cos_I3743 (.Y(N11859), .A0(N11942), .A1(N11964), .B0(N12436));
AND2XL cynw_cm_float_cos_I3744 (.Y(N11992), .A(N11942), .B(N12103));
AO21XL cynw_cm_float_cos_I3745 (.Y(N12129), .A0(N12216), .A1(N12239), .B0(N12078));
AND2XL cynw_cm_float_cos_I3746 (.Y(N12271), .A(N12216), .B(N12381));
AO21XL cynw_cm_float_cos_I3747 (.Y(N12410), .A0(N11863), .A1(N11885), .B0(N12357));
AND2XL cynw_cm_float_cos_I3748 (.Y(N11915), .A(N11863), .B(N12021));
AO21XL cynw_cm_float_cos_I3749 (.Y(N12050), .A0(N12136), .A1(N12159), .B0(N11997));
AND2XL cynw_cm_float_cos_I3750 (.Y(N12190), .A(N12136), .B(N12298));
AO21XL cynw_cm_float_cos_I3751 (.Y(N12329), .A0(N12414), .A1(N12436), .B0(N12275));
AND2XL cynw_cm_float_cos_I3752 (.Y(N11839), .A(N12414), .B(N11942));
AO21XL cynw_cm_float_cos_I3753 (.Y(N11973), .A0(N12054), .A1(N12078), .B0(N11920));
AND2XL cynw_cm_float_cos_I3754 (.Y(N12111), .A(N12054), .B(N12216));
AO21XL cynw_cm_float_cos_I3755 (.Y(N12246), .A0(N12334), .A1(N12357), .B0(N12194));
AND2XL cynw_cm_float_cos_I3756 (.Y(N12390), .A(N12334), .B(N11863));
AO21XL cynw_cm_float_cos_I3757 (.Y(N11892), .A0(N11977), .A1(N11997), .B0(N11843));
AND2XL cynw_cm_float_cos_I3758 (.Y(N12027), .A(N11977), .B(N12136));
AO21XL cynw_cm_float_cos_I3759 (.Y(N12168), .A0(N12250), .A1(N12275), .B0(N12115));
AND2XL cynw_cm_float_cos_I3760 (.Y(N12306), .A(N12250), .B(N12414));
AO21XL cynw_cm_float_cos_I3761 (.Y(N12444), .A0(N11896), .A1(N11920), .B0(N12394));
AND2XL cynw_cm_float_cos_I3762 (.Y(N11950), .A(N11896), .B(N12054));
AO21XL cynw_cm_float_cos_I3763 (.Y(N12086), .A0(N12172), .A1(N12194), .B0(N12031));
AND2XL cynw_cm_float_cos_I3764 (.Y(N12222), .A(N12172), .B(N12334));
AO21XL cynw_cm_float_cos_I3765 (.Y(N12367), .A0(N12448), .A1(N11843), .B0(N12310));
AND2XL cynw_cm_float_cos_I3766 (.Y(N11869), .A(N12448), .B(N11977));
AO21XL cynw_cm_float_cos_I3767 (.Y(N12004), .A0(N12090), .A1(N12115), .B0(N11954));
AND2XL cynw_cm_float_cos_I3768 (.Y(N12144), .A(N12090), .B(N12250));
AO21XL cynw_cm_float_cos_I3769 (.Y(N11957), .A0(N12041), .A1(N12062), .B0(N11906));
AO21XL cynw_cm_float_cos_I3770 (.Y(N12231), .A0(N12318), .A1(N12255), .B0(N12177));
AO21XL cynw_cm_float_cos_I3771 (.Y(N11878), .A0(N11960), .A1(N12092), .B0(N11830));
AO21XL cynw_cm_float_cos_I3772 (.Y(N12151), .A0(N12235), .A1(N12372), .B0(N12100));
AO21XL cynw_cm_float_cos_I3773 (.Y(N12429), .A0(N11881), .A1(N12065), .B0(N12376));
AO21XL cynw_cm_float_cos_I3774 (.Y(N12072), .A0(N12154), .A1(N12345), .B0(N12016));
AO21XL cynw_cm_float_cos_I3775 (.Y(N12268), .A0(N12352), .A1(N11906), .B0(N12212));
AND2XL cynw_cm_float_cos_I3776 (.Y(N12407), .A(N12352), .B(N12041));
AO21XL cynw_cm_float_cos_I3777 (.Y(N11912), .A0(N11992), .A1(N12177), .B0(N11859));
AND2XL cynw_cm_float_cos_I3778 (.Y(N12048), .A(N11992), .B(N12318));
AO21XL cynw_cm_float_cos_I3779 (.Y(N12187), .A0(N12271), .A1(N11830), .B0(N12129));
AND2XL cynw_cm_float_cos_I3780 (.Y(N12326), .A(N12271), .B(N11960));
AO21XL cynw_cm_float_cos_I3781 (.Y(N11837), .A0(N11915), .A1(N12100), .B0(N12410));
AND2XL cynw_cm_float_cos_I3782 (.Y(N11969), .A(N11915), .B(N12235));
AO21XL cynw_cm_float_cos_I3783 (.Y(N12106), .A0(N12190), .A1(N12376), .B0(N12050));
AND2XL cynw_cm_float_cos_I3784 (.Y(N12244), .A(N12190), .B(N11881));
AO21XL cynw_cm_float_cos_I3785 (.Y(N12386), .A0(N11839), .A1(N12016), .B0(N12329));
AND2XL cynw_cm_float_cos_I3786 (.Y(N11889), .A(N11839), .B(N12154));
AO21XL cynw_cm_float_cos_I3787 (.Y(N12024), .A0(N12111), .A1(N12294), .B0(N11973));
AND2XL cynw_cm_float_cos_I3788 (.Y(N12165), .A(N12111), .B(N12432));
AO21XL cynw_cm_float_cos_I3789 (.Y(N12301), .A0(N12390), .A1(N11937), .B0(N12246));
AND2XL cynw_cm_float_cos_I3790 (.Y(N12440), .A(N12390), .B(N12074));
AO21XL cynw_cm_float_cos_I3791 (.Y(N11947), .A0(N12027), .A1(N12212), .B0(N11892));
AND2XL cynw_cm_float_cos_I3792 (.Y(N12083), .A(N12027), .B(N12352));
AO21XL cynw_cm_float_cos_I3793 (.Y(N12219), .A0(N12306), .A1(N11859), .B0(N12168));
AND2XL cynw_cm_float_cos_I3794 (.Y(N12363), .A(N12306), .B(N11992));
AO21XL cynw_cm_float_cos_I3795 (.Y(N11866), .A0(N11950), .A1(N12129), .B0(N12444));
AND2XL cynw_cm_float_cos_I3796 (.Y(N12001), .A(N11950), .B(N12271));
AO21XL cynw_cm_float_cos_I3797 (.Y(N12141), .A0(N12222), .A1(N12410), .B0(N12086));
AND2XL cynw_cm_float_cos_I3798 (.Y(N12280), .A(N12222), .B(N11915));
AO21XL cynw_cm_float_cos_I3799 (.Y(N12417), .A0(N11869), .A1(N12050), .B0(N12367));
AND2XL cynw_cm_float_cos_I3800 (.Y(N11926), .A(N11869), .B(N12190));
AO21XL cynw_cm_float_cos_I3801 (.Y(N12057), .A0(N12144), .A1(N12329), .B0(N12004));
AND2XL cynw_cm_float_cos_I3802 (.Y(N12199), .A(N12144), .B(N11839));
AOI21XL cynw_cm_float_cos_I3803 (.Y(N11930), .A0(N12432), .A1(N11982), .B0(N12294));
AOI21XL cynw_cm_float_cos_I3804 (.Y(N12061), .A0(N12074), .A1(N12261), .B0(N11937));
AO21XL cynw_cm_float_cos_I3805 (.Y(N12323), .A0(N12407), .A1(N12062), .B0(N12268));
AO21XL cynw_cm_float_cos_I3806 (.Y(N11966), .A0(N12048), .A1(N12255), .B0(N11912));
AO21XL cynw_cm_float_cos_I3807 (.Y(N12242), .A0(N12326), .A1(N12092), .B0(N12187));
AO21XL cynw_cm_float_cos_I3808 (.Y(N11887), .A0(N11969), .A1(N12372), .B0(N11837));
AO21XL cynw_cm_float_cos_I3809 (.Y(N12161), .A0(N12244), .A1(N12065), .B0(N12106));
AO21XL cynw_cm_float_cos_I3810 (.Y(N12438), .A0(N11889), .A1(N12345), .B0(N12386));
AO21XL cynw_cm_float_cos_I3811 (.Y(N12080), .A0(N12165), .A1(N11982), .B0(N12024));
AO21XL cynw_cm_float_cos_I3812 (.Y(N12359), .A0(N12440), .A1(N12261), .B0(N12301));
AO21XL cynw_cm_float_cos_I3813 (.Y(N11999), .A0(N12083), .A1(N11957), .B0(N11947));
AO21XL cynw_cm_float_cos_I3814 (.Y(N12277), .A0(N12363), .A1(N12231), .B0(N12219));
AO21XL cynw_cm_float_cos_I3815 (.Y(N11922), .A0(N12001), .A1(N11878), .B0(N11866));
AO21XL cynw_cm_float_cos_I3816 (.Y(N12196), .A0(N12280), .A1(N12151), .B0(N12141));
AO21XL cynw_cm_float_cos_I3817 (.Y(N11846), .A0(N11926), .A1(N12429), .B0(N12417));
AO21XL cynw_cm_float_cos_I3818 (.Y(inst_cellmath__201[49]), .A0(N12199), .A1(N12072), .B0(N12057));
NAND2BXL cynw_cm_float_cos_I3824 (.Y(N11985), .AN(N11827), .B(N11958));
NAND2BXL cynw_cm_float_cos_I3825 (.Y(N12402), .AN(N12099), .B(N12232));
NAND2BXL cynw_cm_float_cos_I3826 (.Y(N12181), .AN(N12374), .B(N11880));
NAND2BXL cynw_cm_float_cos_I3827 (.Y(N11963), .AN(N12014), .B(N12152));
NAND2BXL cynw_cm_float_cos_I3828 (.Y(N12380), .AN(N12293), .B(N12430));
NAND2BXL cynw_cm_float_cos_I3829 (.Y(N12158), .AN(N11935), .B(N12073));
NAND2BXL cynw_cm_float_cos_I3830 (.Y(N11941), .AN(N12210), .B(N12350));
NAND2BXL cynw_cm_float_cos_I3831 (.Y(N12356), .AN(N11858), .B(N11990));
NAND2BXL cynw_cm_float_cos_I3832 (.Y(N12133), .AN(N12127), .B(N12270));
NAND2BXL cynw_cm_float_cos_I3833 (.Y(N11919), .AN(N12408), .B(N11913));
NAND2BXL cynw_cm_float_cos_I3834 (.Y(N12333), .AN(N12049), .B(N12188));
NAND2BXL cynw_cm_float_cos_I3835 (.Y(N12114), .AN(N12327), .B(N11838));
NAND2BXL cynw_cm_float_cos_I3836 (.Y(N11895), .AN(N11971), .B(N12108));
NAND2BXL cynw_cm_float_cos_I3837 (.Y(N12309), .AN(N12245), .B(N12387));
NAND2BXL cynw_cm_float_cos_I3838 (.Y(N12089), .AN(N11890), .B(N12026));
NAND2BXL cynw_cm_float_cos_I3839 (.Y(N11872), .AN(N12166), .B(N12303));
NAND2BXL cynw_cm_float_cos_I3840 (.Y(N12285), .AN(N12442), .B(N11948));
NAND2BXL cynw_cm_float_cos_I3841 (.Y(N12063), .AN(N12084), .B(N12220));
NAND2BXL cynw_cm_float_cos_I3842 (.Y(N11852), .AN(N12364), .B(N11867));
NAND2BXL cynw_cm_float_cos_I3843 (.Y(N12259), .AN(N12002), .B(N12142));
NAND2BXL cynw_cm_float_cos_I3844 (.Y(N12040), .AN(N12281), .B(N12418));
NAND2BXL cynw_cm_float_cos_I3845 (.Y(N11829), .AN(N11928), .B(N12059));
NAND2BXL cynw_cm_float_cos_I3846 (.Y(N12234), .AN(N12200), .B(N12341));
XOR2XL cynw_cm_float_cos_I3852 (.Y(inst_cellmath__201[25]), .A(N12345), .B(N11985));
XOR2XL cynw_cm_float_cos_I3853 (.Y(inst_cellmath__201[26]), .A(N11982), .B(N12402));
XOR2XL cynw_cm_float_cos_I3854 (.Y(inst_cellmath__201[27]), .A(N12261), .B(N12181));
XOR2XL cynw_cm_float_cos_I3855 (.Y(inst_cellmath__201[28]), .A(N11957), .B(N11963));
XOR2XL cynw_cm_float_cos_I3856 (.Y(inst_cellmath__201[29]), .A(N12231), .B(N12380));
XOR2XL cynw_cm_float_cos_I3857 (.Y(inst_cellmath__201[30]), .A(N11878), .B(N12158));
XOR2XL cynw_cm_float_cos_I3858 (.Y(inst_cellmath__201[31]), .A(N12151), .B(N11941));
XOR2XL cynw_cm_float_cos_I3859 (.Y(inst_cellmath__201[32]), .A(N12429), .B(N12356));
XOR2XL cynw_cm_float_cos_I3860 (.Y(inst_cellmath__201[33]), .A(N12072), .B(N12133));
XNOR2X1 cynw_cm_float_cos_I3861 (.Y(inst_cellmath__201[34]), .A(N11930), .B(N11919));
XNOR2X1 cynw_cm_float_cos_I3862 (.Y(inst_cellmath__201[35]), .A(N12061), .B(N12333));
XOR2XL cynw_cm_float_cos_I3863 (.Y(inst_cellmath__201[36]), .A(N12323), .B(N12114));
XOR2XL cynw_cm_float_cos_I3864 (.Y(inst_cellmath__201[37]), .A(N11966), .B(N11895));
XOR2XL cynw_cm_float_cos_I3865 (.Y(inst_cellmath__201[38]), .A(N12242), .B(N12309));
XOR2XL cynw_cm_float_cos_I3866 (.Y(inst_cellmath__201[39]), .A(N11887), .B(N12089));
XOR2XL cynw_cm_float_cos_I3867 (.Y(inst_cellmath__201[40]), .A(N12161), .B(N11872));
XOR2XL cynw_cm_float_cos_I3868 (.Y(inst_cellmath__201[41]), .A(N12438), .B(N12285));
XOR2XL cynw_cm_float_cos_I3869 (.Y(inst_cellmath__201[42]), .A(N12080), .B(N12063));
XOR2XL cynw_cm_float_cos_I3870 (.Y(inst_cellmath__201[43]), .A(N12359), .B(N11852));
XOR2XL cynw_cm_float_cos_I3871 (.Y(inst_cellmath__201[44]), .A(N11999), .B(N12259));
XOR2XL cynw_cm_float_cos_I3872 (.Y(inst_cellmath__201[45]), .A(N12277), .B(N12040));
XOR2XL cynw_cm_float_cos_I3873 (.Y(inst_cellmath__201[46]), .A(N11922), .B(N11829));
XOR2XL cynw_cm_float_cos_I3874 (.Y(inst_cellmath__201[47]), .A(N12196), .B(N12234));
XNOR2X1 cynw_cm_float_cos_I3875 (.Y(inst_cellmath__201[48]), .A(N11846), .B(N12317));
NOR2BX1 cynw_cm_float_cos_I3902 (.Y(inst_cellmath__210[0]), .AN(inst_cellmath__201[25]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3903 (.Y(inst_cellmath__210[1]), .AN(inst_cellmath__201[26]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3904 (.Y(inst_cellmath__210[2]), .AN(inst_cellmath__201[27]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3905 (.Y(inst_cellmath__210[3]), .AN(inst_cellmath__201[28]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3906 (.Y(inst_cellmath__210[4]), .AN(inst_cellmath__201[29]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3907 (.Y(inst_cellmath__210[5]), .AN(inst_cellmath__201[30]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3908 (.Y(inst_cellmath__210[6]), .AN(inst_cellmath__201[31]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3909 (.Y(inst_cellmath__210[7]), .AN(inst_cellmath__201[32]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3910 (.Y(inst_cellmath__210[8]), .AN(inst_cellmath__201[33]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3911 (.Y(inst_cellmath__210[9]), .AN(inst_cellmath__201[34]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3912 (.Y(inst_cellmath__210[10]), .AN(inst_cellmath__201[35]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3913 (.Y(inst_cellmath__210[11]), .AN(inst_cellmath__201[36]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3914 (.Y(inst_cellmath__210[12]), .AN(inst_cellmath__201[37]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3915 (.Y(inst_cellmath__210[13]), .AN(inst_cellmath__201[38]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3916 (.Y(inst_cellmath__210[14]), .AN(inst_cellmath__201[39]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3917 (.Y(inst_cellmath__210[15]), .AN(inst_cellmath__201[40]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3918 (.Y(inst_cellmath__210[16]), .AN(inst_cellmath__201[41]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3919 (.Y(inst_cellmath__210[17]), .AN(inst_cellmath__201[42]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3920 (.Y(inst_cellmath__210[18]), .AN(inst_cellmath__201[43]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3921 (.Y(inst_cellmath__210[19]), .AN(inst_cellmath__201[44]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3922 (.Y(inst_cellmath__210[20]), .AN(inst_cellmath__201[45]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3923 (.Y(inst_cellmath__210[21]), .AN(inst_cellmath__201[46]), .B(inst_cellmath__201[49]));
NOR2BX1 cynw_cm_float_cos_I3924 (.Y(inst_cellmath__210[22]), .AN(inst_cellmath__201[47]), .B(inst_cellmath__201[49]));
OR4X1 inst_cellmath__17_0_I23532 (.Y(N13110), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 inst_cellmath__17_0_I23533 (.Y(N13114), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NOR2XL inst_cellmath__17_0_I3932 (.Y(inst_cellmath__17), .A(N13110), .B(N13114));
NOR2XL andori2bb1_A_I8390 (.Y(N18845), .A(inst_cellmath__42[7]), .B(inst_cellmath__42[6]));
NOR2XL andori2bb1_A_I8391 (.Y(inst_cellmath__46), .A(N18845), .B(inst_cellmath__42[8]));
AOI211XL inst_cellmath__21_0_I3935 (.Y(N13141), .A0(a_exp[2]), .A1(a_exp[1]), .B0(a_exp[3]), .C0(a_exp[4]));
NAND3BXL inst_cellmath__21_0_I3936 (.Y(N13138), .AN(N13141), .B(a_exp[5]), .C(a_exp[6]));
NOR2BX1 inst_cellmath__21_0_I3937 (.Y(inst_cellmath__21), .AN(N13138), .B(a_exp[7]));
OR3XL cynw_cm_float_cos_I3938 (.Y(N494), .A(inst_cellmath__17), .B(inst_cellmath__21), .C(inst_cellmath__46));
NAND2XL inst_cellmath__19_0_I3939 (.Y(N13161), .A(a_exp[7]), .B(a_exp[0]));
AND4XL inst_cellmath__19_0_I23534 (.Y(N13163), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL hyperpropagate_4_1_A_I8392 (.Y(N18854), .A(a_exp[6]), .B(a_exp[5]), .C(N13163));
NOR2XL hyperpropagate_4_1_A_I8393 (.Y(inst_cellmath__19), .A(N13161), .B(N18854));
NOR2XL inst_cellmath__24_0_I3952 (.Y(N13184), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__24_0_I3953 (.Y(N13192), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__24_0_I3954 (.Y(N13203), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__24_0_I3955 (.Y(N13212), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__24_0_I23535 (.Y(N13197), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__24_0_I23536 (.Y(N13206), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__24_0_I23537 (.Y(N13216), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__24_0_I3959 (.Y(N13201), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N13197));
NAND4XL inst_cellmath__24_0_I3961 (.Y(N13195), .A(N13184), .B(N13203), .C(N13192), .D(N13212));
NOR4BX1 inst_cellmath__24_0_I23538 (.Y(inst_cellmath__24), .AN(N13201), .B(N13195), .C(N13206), .D(N13216));
INVXL buf1_A_I8394 (.Y(N18861), .A(inst_cellmath__19));
INVXL buf1_A_I8395 (.Y(inst_cellmath__82), .A(N18861));
AND2XL cynw_cm_float_cos_I23539 (.Y(inst_cellmath__68), .A(inst_cellmath__19), .B(inst_cellmath__24));
OR3XL cynw_cm_float_cos_I3970 (.Y(N741), .A(inst_cellmath__82), .B(inst_cellmath__68), .C(N494));
NAND2XL cynw_cm_float_cos_I8396 (.Y(N18865), .A(inst_cellmath__201[48]), .B(inst_cellmath__61[22]));
INVXL inst_cellmath__211__182__I3972 (.Y(N13336), .A(inst_cellmath__210[22]));
INVXL inst_cellmath__211__182__I3973 (.Y(N13278), .A(inst_cellmath__210[0]));
INVXL inst_cellmath__211__182__I3974 (.Y(N13314), .A(inst_cellmath__210[2]));
OAI21XL inst_cellmath__211__182__I3975 (.Y(N13331), .A0(inst_cellmath__210[1]), .A1(N13278), .B0(N13314));
OR2XL inst_cellmath__211__182__I3976 (.Y(N13335), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[1]));
NOR2BX1 inst_cellmath__211__182__I3977 (.Y(N13322), .AN(inst_cellmath__210[3]), .B(inst_cellmath__210[4]));
INVXL inst_cellmath__211__182__I3978 (.Y(N13340), .A(inst_cellmath__210[6]));
OAI21XL inst_cellmath__211__182__I3979 (.Y(N13275), .A0(inst_cellmath__210[5]), .A1(N13322), .B0(N13340));
NOR2XL inst_cellmath__211__182__I3980 (.Y(N13293), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[3]));
NOR2XL inst_cellmath__211__182__I3981 (.Y(N13309), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[5]));
NOR2BX1 inst_cellmath__211__182__I3982 (.Y(N13347), .AN(inst_cellmath__210[7]), .B(inst_cellmath__210[8]));
INVXL inst_cellmath__211__182__I3983 (.Y(N13281), .A(inst_cellmath__210[10]));
OAI21XL inst_cellmath__211__182__I3984 (.Y(N13300), .A0(inst_cellmath__210[9]), .A1(N13347), .B0(N13281));
NOR2XL inst_cellmath__211__182__I3985 (.Y(N13318), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[7]));
NOR2XL inst_cellmath__211__182__I3986 (.Y(N13337), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[9]));
NOR2BX1 inst_cellmath__211__182__I3987 (.Y(N13290), .AN(inst_cellmath__210[11]), .B(inst_cellmath__210[12]));
INVXL inst_cellmath__211__182__I3988 (.Y(N13306), .A(inst_cellmath__210[14]));
OAI21XL inst_cellmath__211__182__I3989 (.Y(N13326), .A0(inst_cellmath__210[13]), .A1(N13290), .B0(N13306));
NOR2XL inst_cellmath__211__182__I3990 (.Y(N13345), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[11]));
NOR2XL inst_cellmath__211__182__I3991 (.Y(N13279), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[13]));
NOR2BX1 inst_cellmath__211__182__I3992 (.Y(N13315), .AN(inst_cellmath__210[15]), .B(inst_cellmath__210[16]));
INVXL inst_cellmath__211__182__I3993 (.Y(N13333), .A(inst_cellmath__210[18]));
OAI21XL inst_cellmath__211__182__I3994 (.Y(N13270), .A0(inst_cellmath__210[17]), .A1(N13315), .B0(N13333));
NOR2XL inst_cellmath__211__182__I3995 (.Y(N13286), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[15]));
NOR2XL inst_cellmath__211__182__I3996 (.Y(N13303), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[17]));
NOR2BX1 inst_cellmath__211__182__I3997 (.Y(N13342), .AN(inst_cellmath__210[19]), .B(inst_cellmath__210[20]));
OAI21XL inst_cellmath__211__182__I3998 (.Y(N13296), .A0(inst_cellmath__210[21]), .A1(N13342), .B0(N13336));
NOR2XL inst_cellmath__211__182__I3999 (.Y(N13311), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[19]));
NOR2XL inst_cellmath__211__182__I4000 (.Y(N13329), .A(inst_cellmath__210[22]), .B(inst_cellmath__210[21]));
INVXL inst_cellmath__211__182__I4001 (.Y(N13287), .A(N13309));
AOI21XL inst_cellmath__211__182__I4002 (.Y(N13305), .A0(N13293), .A1(N13335), .B0(N13287));
NAND2XL inst_cellmath__211__182__I4003 (.Y(N13343), .A(N13309), .B(N13293));
NAND2BXL inst_cellmath__211__182__I4004 (.Y(N13297), .AN(N13318), .B(N13337));
INVXL inst_cellmath__211__182__I4005 (.Y(N13313), .A(N13279));
AOI21XL inst_cellmath__211__182__I4006 (.Y(N13330), .A0(N13345), .A1(N13297), .B0(N13313));
NAND2XL inst_cellmath__211__182__I4007 (.Y(N13349), .A(N13337), .B(N13318));
NAND2XL inst_cellmath__211__182__I4008 (.Y(N13284), .A(N13279), .B(N13345));
NAND2BXL inst_cellmath__211__182__I4009 (.Y(N13321), .AN(N13286), .B(N13303));
NAND2XL inst_cellmath__211__182__I4010 (.Y(N13292), .A(N13303), .B(N13286));
NAND2XL inst_cellmath__211__182__I4011 (.Y(N13308), .A(N13329), .B(N13311));
INVXL inst_cellmath__211__182__I4012 (.Y(N13289), .A(N13343));
INVXL inst_cellmath__211__182__I4013 (.Y(N13325), .A(N13284));
OAI21XL inst_cellmath__211__182__I4014 (.Y(N13344), .A0(N13349), .A1(N13289), .B0(N13325));
NOR2XL inst_cellmath__211__182__I4015 (.Y(N13294), .A(N13284), .B(N13349));
NAND2BXL inst_cellmath__211__182__I4016 (.Y(N13285), .AN(N13308), .B(N13292));
OR2XL inst_cellmath__211__182__I4017 (.Y(N13324), .A(N13308), .B(N13292));
OR2XL inst_cellmath__211__182__I4018 (.Y(N551), .A(N13324), .B(N13294));
OAI21XL inst_cellmath__211__182__I4020 (.Y(N550), .A0(N13324), .A1(N13344), .B0(N13285));
AOI21XL inst_cellmath__211__182__I4021 (.Y(N13277), .A0(N13294), .A1(N13305), .B0(N13330));
OAI2BB1X1 inst_cellmath__211__182__I4022 (.Y(N13312), .A0N(N13311), .A1N(N13321), .B0(N13329));
OAI21XL inst_cellmath__211__182__I4023 (.Y(N549), .A0(N13324), .A1(N13277), .B0(N13312));
OAI21XL inst_cellmath__211__182__I4024 (.Y(N13317), .A0(N13343), .A1(N13331), .B0(N13275));
OAI21XL inst_cellmath__211__182__I4025 (.Y(N13272), .A0(N13284), .A1(N13300), .B0(N13326));
AOI21XL inst_cellmath__211__182__I4026 (.Y(N13298), .A0(N13294), .A1(N13317), .B0(N13272));
OA21X1 inst_cellmath__211__182__I4027 (.Y(N13332), .A0(N13270), .A1(N13308), .B0(N13296));
OAI21XL inst_cellmath__211__182__I4028 (.Y(N548), .A0(N13324), .A1(N13298), .B0(N13332));
INVXL inst_cellmath__215_0_I4029 (.Y(inst_cellmath__215[0]), .A(N548));
NAND2XL inst_cellmath__215_0_I4030 (.Y(N13410), .A(N549), .B(N548));
NAND3XL inst_cellmath__215_0_I4031 (.Y(N13408), .A(N550), .B(N549), .C(N548));
NAND2BXL inst_cellmath__215_0_I4032 (.Y(N13413), .AN(N551), .B(N13408));
XOR2XL inst_cellmath__215_0_I4035 (.Y(inst_cellmath__215[3]), .A(N13408), .B(N551));
INVXL inst_cellmath__220__188__I4037 (.Y(N13539), .A(inst_cellmath__215[0]));
AND2XL inst_cellmath__220__188__I4038 (.Y(N13577), .A(N13539), .B(inst_cellmath__210[0]));
MX2XL inst_cellmath__220__188__I4039 (.Y(N13493), .A(inst_cellmath__210[0]), .B(inst_cellmath__210[1]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4040 (.Y(N13527), .A(inst_cellmath__210[1]), .B(inst_cellmath__210[2]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4041 (.Y(N13561), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[3]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4042 (.Y(N13441), .A(inst_cellmath__210[3]), .B(inst_cellmath__210[4]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4043 (.Y(N13472), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[5]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4044 (.Y(N13509), .A(inst_cellmath__210[5]), .B(inst_cellmath__210[6]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4045 (.Y(N13542), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[7]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4046 (.Y(N13573), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4047 (.Y(N13456), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[9]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4048 (.Y(N13486), .A(inst_cellmath__210[9]), .B(inst_cellmath__210[10]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4049 (.Y(N13521), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[11]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4050 (.Y(N13555), .A(inst_cellmath__210[11]), .B(inst_cellmath__210[12]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4051 (.Y(N13435), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[13]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4052 (.Y(N13465), .A(inst_cellmath__210[13]), .B(inst_cellmath__210[14]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4053 (.Y(N13503), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[15]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4054 (.Y(N13536), .A(inst_cellmath__210[15]), .B(inst_cellmath__210[16]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4055 (.Y(N13567), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[17]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4056 (.Y(N13450), .A(inst_cellmath__210[17]), .B(inst_cellmath__210[18]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4057 (.Y(N13479), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[19]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4058 (.Y(N13515), .A(inst_cellmath__210[19]), .B(inst_cellmath__210[20]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4059 (.Y(N13550), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[21]), .S0(N13539));
MX2XL inst_cellmath__220__188__I4060 (.Y(N13430), .A(inst_cellmath__210[21]), .B(inst_cellmath__210[22]), .S0(N13539));
XOR2XL inst_cellmath__220__188__I8352 (.Y(N13532), .A(inst_cellmath__215[0]), .B(N549));
INVXL inst_cellmath__220__188__I4062 (.Y(N13547), .A(N13532));
NAND2XL inst_cellmath__220__188__I4063 (.Y(N13445), .A(N13577), .B(N13532));
NAND2XL inst_cellmath__220__188__I4064 (.Y(N13512), .A(N13493), .B(N13532));
AOI22XL inst_cellmath__220__188__I4065 (.Y(N13576), .A0(N13547), .A1(N13577), .B0(N13527), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4066 (.Y(N13459), .A0(N13547), .A1(N13493), .B0(N13561), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4067 (.Y(N13492), .A0(N13547), .A1(N13527), .B0(N13441), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4068 (.Y(N13525), .A0(N13547), .A1(N13561), .B0(N13472), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4069 (.Y(N13559), .A0(N13547), .A1(N13441), .B0(N13509), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4070 (.Y(N13440), .A0(N13547), .A1(N13472), .B0(N13542), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4071 (.Y(N13471), .A0(N13547), .A1(N13509), .B0(N13573), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4072 (.Y(N13508), .A0(N13547), .A1(N13542), .B0(N13456), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4073 (.Y(N13541), .A0(N13547), .A1(N13573), .B0(N13486), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4074 (.Y(N13572), .A0(N13547), .A1(N13456), .B0(N13521), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4075 (.Y(N13455), .A0(N13547), .A1(N13486), .B0(N13555), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4076 (.Y(N13485), .A0(N13547), .A1(N13521), .B0(N13435), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4077 (.Y(N13520), .A0(N13547), .A1(N13555), .B0(N13465), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4078 (.Y(N13554), .A0(N13547), .A1(N13435), .B0(N13503), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4079 (.Y(N13434), .A0(N13547), .A1(N13465), .B0(N13536), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4080 (.Y(N13464), .A0(N13547), .A1(N13503), .B0(N13567), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4081 (.Y(N13501), .A0(N13547), .A1(N13536), .B0(N13450), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4082 (.Y(N13534), .A0(N13547), .A1(N13567), .B0(N13479), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4083 (.Y(N13566), .A0(N13547), .A1(N13450), .B0(N13515), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4084 (.Y(N13449), .A0(N13547), .A1(N13479), .B0(N13550), .B1(N13532));
AOI22XL inst_cellmath__220__188__I4085 (.Y(N13478), .A0(N13547), .A1(N13515), .B0(N13430), .B1(N13532));
XOR2XL inst_cellmath__220__188__I8353 (.Y(N13487), .A(N13410), .B(N550));
INVXL inst_cellmath__220__188__I4087 (.Y(N13504), .A(N13487));
NOR2XL inst_cellmath__220__188__I4088 (.Y(N13498), .A(N13504), .B(N13445));
NOR2XL inst_cellmath__220__188__I4089 (.Y(N13444), .A(N13504), .B(N13512));
NOR2XL inst_cellmath__220__188__I4090 (.Y(N13546), .A(N13504), .B(N13576));
NOR2XL inst_cellmath__220__188__I4091 (.Y(N13491), .A(N13504), .B(N13459));
AOI22XL inst_cellmath__220__188__I4092 (.Y(N13439), .A0(N13487), .A1(N13492), .B0(N13445), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4093 (.Y(N13470), .A0(N13487), .A1(N13525), .B0(N13512), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4094 (.Y(N13507), .A0(N13487), .A1(N13559), .B0(N13576), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4095 (.Y(N13540), .A0(N13487), .A1(N13440), .B0(N13459), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4096 (.Y(N13571), .A0(N13487), .A1(N13471), .B0(N13492), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4097 (.Y(N13454), .A0(N13487), .A1(N13508), .B0(N13525), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4098 (.Y(N13484), .A0(N13487), .A1(N13541), .B0(N13559), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4099 (.Y(N13519), .A0(N13487), .A1(N13572), .B0(N13440), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4100 (.Y(N13553), .A0(N13487), .A1(N13455), .B0(N13471), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4101 (.Y(N13433), .A0(N13487), .A1(N13485), .B0(N13508), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4102 (.Y(N13463), .A0(N13487), .A1(N13520), .B0(N13541), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4103 (.Y(N13500), .A0(N13487), .A1(N13554), .B0(N13572), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4104 (.Y(N13533), .A0(N13487), .A1(N13434), .B0(N13455), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4105 (.Y(N13565), .A0(N13487), .A1(N13464), .B0(N13485), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4106 (.Y(N13448), .A0(N13487), .A1(N13501), .B0(N13520), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4107 (.Y(N13477), .A0(N13487), .A1(N13534), .B0(N13554), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4108 (.Y(N13514), .A0(N13487), .A1(N13566), .B0(N13434), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4109 (.Y(N13548), .A0(N13487), .A1(N13449), .B0(N13464), .B1(N13504));
AOI22XL inst_cellmath__220__188__I4110 (.Y(N13428), .A0(N13487), .A1(N13478), .B0(N13501), .B1(N13504));
INVXL inst_cellmath__220__188__I4111 (.Y(N13489), .A(inst_cellmath__215[3]));
NAND2XL inst_cellmath__220__188__I4112 (.Y(N13447), .A(N13498), .B(N13489));
NAND2XL inst_cellmath__220__188__I4113 (.Y(N13513), .A(N13444), .B(N13489));
NAND2XL inst_cellmath__220__188__I4114 (.Y(N13578), .A(N13546), .B(N13489));
NAND2XL inst_cellmath__220__188__I4115 (.Y(N13494), .A(N13491), .B(N13489));
NAND2XL inst_cellmath__220__188__I4116 (.Y(N13560), .A(N13439), .B(N13489));
NAND2XL inst_cellmath__220__188__I4117 (.Y(N13473), .A(N13470), .B(N13489));
NAND2XL inst_cellmath__220__188__I4118 (.Y(N13543), .A(N13507), .B(N13489));
AOI22XL inst_cellmath__220__188__I4119 (.Y(N13522), .A0(inst_cellmath__215[3]), .A1(N13498), .B0(N13571), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4120 (.Y(N13556), .A0(inst_cellmath__215[3]), .A1(N13444), .B0(N13454), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4121 (.Y(N13436), .A0(inst_cellmath__215[3]), .A1(N13546), .B0(N13484), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4122 (.Y(N13466), .A0(inst_cellmath__215[3]), .A1(N13491), .B0(N13519), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4123 (.Y(N13502), .A0(inst_cellmath__215[3]), .A1(N13439), .B0(N13553), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4124 (.Y(N13535), .A0(inst_cellmath__215[3]), .A1(N13470), .B0(N13433), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4125 (.Y(N13568), .A0(inst_cellmath__215[3]), .A1(N13507), .B0(N13463), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4126 (.Y(N13451), .A0(inst_cellmath__215[3]), .A1(N13540), .B0(N13500), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4127 (.Y(N13480), .A0(inst_cellmath__215[3]), .A1(N13571), .B0(N13533), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4128 (.Y(N13516), .A0(inst_cellmath__215[3]), .A1(N13454), .B0(N13565), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4129 (.Y(N13549), .A0(inst_cellmath__215[3]), .A1(N13484), .B0(N13448), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4130 (.Y(N13429), .A0(inst_cellmath__215[3]), .A1(N13519), .B0(N13477), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4131 (.Y(N13460), .A0(inst_cellmath__215[3]), .A1(N13553), .B0(N13514), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4132 (.Y(N13496), .A0(inst_cellmath__215[3]), .A1(N13433), .B0(N13548), .B1(N13489));
AOI22XL inst_cellmath__220__188__I4133 (.Y(N13529), .A0(inst_cellmath__215[3]), .A1(N13463), .B0(N13428), .B1(N13489));
XNOR2X1 inst_cellmath__220__188__I8354 (.Y(N13469), .A(N13413), .B(N13324));
INVXL inst_cellmath__220__188__I4135 (.Y(N13483), .A(N13469));
AOI22XL inst_cellmath__220__188__I4153 (.Y(N677), .A0(N13469), .A1(N13480), .B0(N13447), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4154 (.Y(N678), .A0(N13469), .A1(N13516), .B0(N13513), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4155 (.Y(N679), .A0(N13469), .A1(N13549), .B0(N13578), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4156 (.Y(N680), .A0(N13469), .A1(N13429), .B0(N13494), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4157 (.Y(N681), .A0(N13469), .A1(N13460), .B0(N13560), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4158 (.Y(N682), .A0(N13469), .A1(N13496), .B0(N13473), .B1(N13483));
AOI22XL inst_cellmath__220__188__I4159 (.Y(N683), .A0(N13469), .A1(N13529), .B0(N13543), .B1(N13483));
OR2XL inst_cellmath__220_2WWMM_I23540 (.Y(N13757), .A(inst_cellmath__201[49]), .B(N18865));
NAND2BXL inst_cellmath__220_2WWMM_I4166 (.Y(N709), .AN(N13539), .B(N13757));
NAND2BXL inst_cellmath__220_2WWMM_I4167 (.Y(N710), .AN(N13532), .B(N13757));
NAND2BXL inst_cellmath__220_2WWMM_I4168 (.Y(N711), .AN(N13487), .B(N13757));
NAND2BXL inst_cellmath__220_2WWMM_I4169 (.Y(N712), .AN(N13489), .B(N13757));
NAND2BXL inst_cellmath__220_2WWMM_I4170 (.Y(N713), .AN(N13469), .B(N13757));
NOR3BXL inst_cellmath__220_2WWMM_I8356 (.Y(N717), .AN(N13757), .B(N13483), .C(N13447));
NOR3BXL inst_cellmath__220_2WWMM_I8357 (.Y(N718), .AN(N13757), .B(N13483), .C(N13513));
NOR3BXL inst_cellmath__220_2WWMM_I8358 (.Y(N719), .AN(N13757), .B(N13483), .C(N13578));
NOR3BXL inst_cellmath__220_2WWMM_I8359 (.Y(N720), .AN(N13757), .B(N13483), .C(N13494));
NOR3BXL inst_cellmath__220_2WWMM_I8360 (.Y(N721), .AN(N13757), .B(N13483), .C(N13560));
NOR3BXL inst_cellmath__220_2WWMM_I8361 (.Y(N722), .AN(N13757), .B(N13483), .C(N13473));
NOR3BXL inst_cellmath__220_2WWMM_I8362 (.Y(N723), .AN(N13757), .B(N13483), .C(N13543));
NAND3XL hyperpropagate_4_1_A_I8398 (.Y(N18874), .A(N13540), .B(N13757), .C(N13489));
NOR2XL hyperpropagate_4_1_A_I8399 (.Y(N724), .A(N13483), .B(N18874));
NOR3BXL inst_cellmath__220_2WWMM_I8364 (.Y(N725), .AN(N13757), .B(N13483), .C(N13522));
NOR3BXL inst_cellmath__220_2WWMM_I8365 (.Y(N726), .AN(N13757), .B(N13483), .C(N13556));
NOR3BXL inst_cellmath__220_2WWMM_I8366 (.Y(N727), .AN(N13757), .B(N13483), .C(N13436));
NOR3BXL inst_cellmath__220_2WWMM_I8367 (.Y(N728), .AN(N13757), .B(N13483), .C(N13466));
NOR3BXL inst_cellmath__220_2WWMM_I8368 (.Y(N729), .AN(N13757), .B(N13483), .C(N13502));
NOR3BXL inst_cellmath__220_2WWMM_I8369 (.Y(N730), .AN(N13757), .B(N13483), .C(N13535));
NOR3BXL inst_cellmath__220_2WWMM_I8370 (.Y(N731), .AN(N13757), .B(N13483), .C(N13568));
NOR3BXL inst_cellmath__220_2WWMM_I8371 (.Y(N732), .AN(N13757), .B(N13483), .C(N13451));
AND2XL inst_cellmath__220_2WWMM_I4189 (.Y(N733), .A(N13757), .B(N677));
AND2XL inst_cellmath__220_2WWMM_I4190 (.Y(N734), .A(N13757), .B(N678));
AND2XL inst_cellmath__220_2WWMM_I4191 (.Y(N735), .A(N13757), .B(N679));
AND2XL inst_cellmath__220_2WWMM_I4192 (.Y(N736), .A(N13757), .B(N680));
AND2XL inst_cellmath__220_2WWMM_I4193 (.Y(N737), .A(N13757), .B(N681));
AND2XL inst_cellmath__220_2WWMM_I4194 (.Y(N738), .A(N13757), .B(N682));
AND2XL inst_cellmath__220_2WWMM_I4195 (.Y(N739), .A(N13757), .B(N683));
NOR2XL inst_cellmath__223__199__I4213 (.Y(N13872), .A(inst_cellmath__42[6]), .B(inst_cellmath__82));
NOR4BBX1 inst_cellmath__223__199__I8372 (.Y(x[31]), .AN(N13872), .BN(N493), .C(inst_cellmath__42[8]), .D(inst_cellmath__42[7]));
OR2XL cynw_cm_float_cos_I4215 (.Y(N585), .A(inst_cellmath__68), .B(N494));
NAND2BXL cynw_cm_float_cos_I4216 (.Y(N595), .AN(inst_cellmath__82), .B(N585));
NAND2BXL cynw_cm_float_cos_I4217 (.Y(N594), .AN(inst_cellmath__82), .B(inst_cellmath__68));
INVXL inst_cellmath__228_0_I4218 (.Y(N13910), .A(N741));
INVXL inst_cellmath__228_0_I4219 (.Y(N13897), .A(N13910));
MX2XL inst_cellmath__228_0_I4220 (.Y(x[23]), .A(N709), .B(N594), .S0(N13897));
MX2XL inst_cellmath__228_0_I4221 (.Y(x[24]), .A(N710), .B(N594), .S0(N13897));
MX2XL inst_cellmath__228_0_I4222 (.Y(x[25]), .A(N711), .B(N594), .S0(N13897));
MX2XL inst_cellmath__228_0_I4223 (.Y(x[26]), .A(N712), .B(N594), .S0(N13897));
MX2XL inst_cellmath__228_0_I4224 (.Y(x[27]), .A(N713), .B(N594), .S0(N13897));
NAND2BXL inst_cellmath__228_0_I4225 (.Y(x[28]), .AN(N594), .B(N13897));
AND2XL inst_cellmath__228_0_I4227 (.Y(x[30]), .A(N13897), .B(N595));
MX2XL inst_cellmath__231_0_I4228 (.Y(x[0]), .A(N717), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4229 (.Y(x[1]), .A(N718), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4230 (.Y(x[2]), .A(N719), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4231 (.Y(x[3]), .A(N720), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4232 (.Y(x[4]), .A(N721), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4233 (.Y(x[5]), .A(N722), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4234 (.Y(x[6]), .A(N723), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4235 (.Y(x[7]), .A(N724), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4236 (.Y(x[8]), .A(N725), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4237 (.Y(x[9]), .A(N726), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4238 (.Y(x[10]), .A(N727), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4239 (.Y(x[11]), .A(N728), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4240 (.Y(x[12]), .A(N729), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4241 (.Y(x[13]), .A(N730), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4242 (.Y(x[14]), .A(N731), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4243 (.Y(x[15]), .A(N732), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4244 (.Y(x[16]), .A(N733), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4245 (.Y(x[17]), .A(N734), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4246 (.Y(x[18]), .A(N735), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4247 (.Y(x[19]), .A(N736), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4248 (.Y(x[20]), .A(N737), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4249 (.Y(x[21]), .A(N738), .B(inst_cellmath__82), .S0(N741));
MX2XL inst_cellmath__231_0_I4250 (.Y(x[22]), .A(N739), .B(inst_cellmath__82), .S0(N741));
assign inst_cellmath__42[0] = 1'B0;
assign inst_cellmath__42[2] = 1'B0;
assign inst_cellmath__42[3] = 1'B0;
assign inst_cellmath__42[5] = 1'B0;
assign inst_cellmath__61[0] = 1'B0;
assign inst_cellmath__61[16] = 1'B0;
assign inst_cellmath__61[19] = 1'B0;
assign inst_cellmath__61[20] = 1'B0;
assign inst_cellmath__61[21] = 1'B0;
assign inst_cellmath__195[29] = 1'B0;
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__198[0] = 1'B0;
assign inst_cellmath__198[1] = 1'B0;
assign inst_cellmath__198[2] = 1'B0;
assign inst_cellmath__198[3] = 1'B0;
assign inst_cellmath__198[4] = 1'B0;
assign inst_cellmath__198[5] = 1'B0;
assign inst_cellmath__198[6] = 1'B0;
assign inst_cellmath__198[7] = 1'B0;
assign inst_cellmath__198[8] = 1'B0;
assign inst_cellmath__198[9] = 1'B0;
assign inst_cellmath__198[10] = 1'B0;
assign inst_cellmath__198[11] = 1'B0;
assign inst_cellmath__198[12] = 1'B0;
assign inst_cellmath__198[13] = 1'B0;
assign inst_cellmath__198[14] = 1'B0;
assign inst_cellmath__198[15] = 1'B0;
assign inst_cellmath__198[16] = 1'B0;
assign inst_cellmath__198[17] = 1'B0;
assign inst_cellmath__201[0] = 1'B0;
assign inst_cellmath__201[1] = 1'B0;
assign inst_cellmath__201[2] = 1'B0;
assign inst_cellmath__201[3] = 1'B0;
assign inst_cellmath__201[4] = 1'B0;
assign inst_cellmath__201[5] = 1'B0;
assign inst_cellmath__201[6] = 1'B0;
assign inst_cellmath__201[7] = 1'B0;
assign inst_cellmath__201[8] = 1'B0;
assign inst_cellmath__201[9] = 1'B0;
assign inst_cellmath__201[10] = 1'B0;
assign inst_cellmath__201[11] = 1'B0;
assign inst_cellmath__201[12] = 1'B0;
assign inst_cellmath__201[13] = 1'B0;
assign inst_cellmath__201[14] = 1'B0;
assign inst_cellmath__201[15] = 1'B0;
assign inst_cellmath__201[16] = 1'B0;
assign inst_cellmath__201[17] = 1'B0;
assign inst_cellmath__201[18] = 1'B0;
assign inst_cellmath__201[19] = 1'B0;
assign inst_cellmath__201[20] = 1'B0;
assign inst_cellmath__201[21] = 1'B0;
assign inst_cellmath__201[22] = 1'B0;
assign inst_cellmath__201[23] = 1'B0;
assign inst_cellmath__201[24] = 1'B0;
assign inst_cellmath__203__W0[0] = 1'B0;
assign inst_cellmath__203__W0[43] = 1'B1;
assign inst_cellmath__203__W0[44] = 1'B1;
assign inst_cellmath__203__W0[45] = 1'B1;
assign inst_cellmath__203__W0[46] = 1'B1;
assign inst_cellmath__203__W1[0] = 1'B0;
assign inst_cellmath__203__W1[43] = 1'B0;
assign inst_cellmath__203__W1[44] = 1'B0;
assign inst_cellmath__203__W1[45] = 1'B0;
assign inst_cellmath__203__W1[46] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign inst_cellmath__215[1] = 1'B0;
assign inst_cellmath__215[2] = 1'B0;
assign inst_cellmath__215[4] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  v7PyTw7aqBw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



