/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:24:33 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46;
wire [22:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874,
	DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297;
wire N18241,N18245,N18402,N18406,N19158,N19431,N19751 
	,N19755,N20260,N20265,N20270,N20275,N20280,N20285,N20290 
	,N20295,N20355,N20370,N20382,N20609,N20613,N20621,N20625 
	,N20628,N20632,N20654,N20872,N20876,N20886,N20890,N20899 
	,N20903,N20912,N20916,N21060,N21064,N21306,N21310,N21559 
	,N21570,N21574,N21818,N21831,N21833,N21853,N21863,N21873 
	,N21883,N21893,N21903,N21913,N21923,N21933,N21943,N21953 
	,N21963,N21973,N21983,N21993,N21997,N22003,N22005,N22007 
	,N22034,N22040,N22048,N22056,N22064,N22066,N22072,N22080 
	,N22082,N22091,N22097,N22101,N22105,N22109,N22113,N22117 
	,N22121,N22123,N22125,N22129,N22131,N22133,N22137,N22139 
	,N22141,N22145,N22147,N22149,N22153,N22155,N22157,N22194 
	,N22199,N22201,N22203,N22205,N22209,N22211,N22213,N22217 
	,N22219,N22221,N22225,N22227,N22229,N22233,N22235,N22237 
	,N22241,N22243,N22245,N22249,N22251,N22253,N22258,N22260 
	,N22268,N22270,N22278,N22286,N22288,N22290,N22294,N22296 
	,N22306,N22310,N22314,N22316,N22318,N22322,N22324,N22326 
	,N22678,N22680,N22961,N22962,N22963,N22964,N22965,N22966 
	,N22968,N22969,N22971;
reg x_reg_22__retimed_I12950_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12950_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250;
	end
assign N22680 = x_reg_22__retimed_I12950_QOUT;
reg x_reg_22__retimed_I12949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12949_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090;
	end
assign N22678 = x_reg_22__retimed_I12949_QOUT;
reg x_reg_22__retimed_I12809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12809_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253;
	end
assign N22326 = x_reg_22__retimed_I12809_QOUT;
reg x_reg_22__retimed_I12808_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12808_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035;
	end
assign N22324 = x_reg_22__retimed_I12808_QOUT;
reg x_reg_22__retimed_I12807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12807_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214;
	end
assign N22322 = x_reg_22__retimed_I12807_QOUT;
reg x_reg_22__retimed_I12806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12806_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673;
	end
assign N22318 = x_reg_22__retimed_I12806_QOUT;
reg x_reg_22__retimed_I12805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12805_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176;
	end
assign N22316 = x_reg_22__retimed_I12805_QOUT;
reg x_reg_22__retimed_I12804_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12804_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633;
	end
assign N22314 = x_reg_22__retimed_I12804_QOUT;
reg x_reg_22__retimed_I12803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12803_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017;
	end
assign N22310 = x_reg_22__retimed_I12803_QOUT;
reg x_reg_22__retimed_I12801_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12801_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999;
	end
assign N22306 = x_reg_22__retimed_I12801_QOUT;
reg x_reg_22__retimed_I12798_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12798_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[14];
	end
assign N22296 = x_reg_22__retimed_I12798_QOUT;
reg x_reg_22__retimed_I12797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12797_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[14];
	end
assign N22294 = x_reg_22__retimed_I12797_QOUT;
reg x_reg_22__retimed_I12796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12796_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642;
	end
assign N22290 = x_reg_22__retimed_I12796_QOUT;
reg x_reg_22__retimed_I12795_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12795_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873;
	end
assign N22288 = x_reg_22__retimed_I12795_QOUT;
reg x_reg_22__retimed_I12794_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12794_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829;
	end
assign N22286 = x_reg_22__retimed_I12794_QOUT;
reg x_reg_22__retimed_I12792_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12792_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[0];
	end
assign N22278 = x_reg_22__retimed_I12792_QOUT;
reg x_reg_22__retimed_I12790_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12790_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005;
	end
assign N22270 = x_reg_22__retimed_I12790_QOUT;
reg x_reg_22__retimed_I12789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12789_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052;
	end
assign N22268 = x_reg_22__retimed_I12789_QOUT;
reg x_reg_22__retimed_I12787_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12787_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402;
	end
assign N22260 = x_reg_22__retimed_I12787_QOUT;
reg x_reg_22__retimed_I12786_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12786_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205;
	end
assign N22258 = x_reg_22__retimed_I12786_QOUT;
reg x_reg_22__retimed_I12785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12785_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143;
	end
assign N22253 = x_reg_22__retimed_I12785_QOUT;
reg x_reg_22__retimed_I12784_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12784_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720;
	end
assign N22251 = x_reg_22__retimed_I12784_QOUT;
reg x_reg_22__retimed_I12783_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12783_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117;
	end
assign N22249 = x_reg_22__retimed_I12783_QOUT;
reg x_reg_22__retimed_I12782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12782_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597;
	end
assign N22245 = x_reg_22__retimed_I12782_QOUT;
reg x_reg_22__retimed_I12781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12781_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140;
	end
assign N22243 = x_reg_22__retimed_I12781_QOUT;
reg x_reg_22__retimed_I12780_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12780_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835;
	end
assign N22241 = x_reg_22__retimed_I12780_QOUT;
reg x_reg_22__retimed_I12779_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12779_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098;
	end
assign N22237 = x_reg_22__retimed_I12779_QOUT;
reg x_reg_22__retimed_I12778_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12778_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073;
	end
assign N22235 = x_reg_22__retimed_I12778_QOUT;
reg x_reg_22__retimed_I12777_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12777_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592;
	end
assign N22233 = x_reg_22__retimed_I12777_QOUT;
reg x_reg_22__retimed_I12776_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12776_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559;
	end
assign N22229 = x_reg_22__retimed_I12776_QOUT;
reg x_reg_22__retimed_I12775_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12775_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130;
	end
assign N22227 = x_reg_22__retimed_I12775_QOUT;
reg x_reg_22__retimed_I12774_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12774_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800;
	end
assign N22225 = x_reg_22__retimed_I12774_QOUT;
reg x_reg_22__retimed_I12773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12773_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257;
	end
assign N22221 = x_reg_22__retimed_I12773_QOUT;
reg x_reg_22__retimed_I12772_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12772_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827;
	end
assign N22219 = x_reg_22__retimed_I12772_QOUT;
reg x_reg_22__retimed_I12771_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12771_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217;
	end
assign N22217 = x_reg_22__retimed_I12771_QOUT;
reg x_reg_22__retimed_I12770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12770_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588;
	end
assign N22213 = x_reg_22__retimed_I12770_QOUT;
reg x_reg_22__retimed_I12769_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12769_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862;
	end
assign N22211 = x_reg_22__retimed_I12769_QOUT;
reg x_reg_22__retimed_I12768_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12768_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521;
	end
assign N22209 = x_reg_22__retimed_I12768_QOUT;
reg x_reg_22__retimed_I12767_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12767_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391;
	end
assign N22205 = x_reg_22__retimed_I12767_QOUT;
reg x_reg_22__retimed_I12766_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12766_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12];
	end
assign N22203 = x_reg_22__retimed_I12766_QOUT;
reg x_reg_22__retimed_I12765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12765_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12];
	end
assign N22201 = x_reg_22__retimed_I12765_QOUT;
reg x_reg_22__retimed_I12764_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12764_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134;
	end
assign N22199 = x_reg_22__retimed_I12764_QOUT;
reg x_reg_22__retimed_I12762_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12762_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893;
	end
assign N22194 = x_reg_22__retimed_I12762_QOUT;
reg x_reg_22__retimed_I12748_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12748_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629;
	end
assign N22157 = x_reg_22__retimed_I12748_QOUT;
reg x_reg_22__retimed_I12747_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12747_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320;
	end
assign N22155 = x_reg_22__retimed_I12747_QOUT;
reg x_reg_22__retimed_I12746_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12746_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578;
	end
assign N22153 = x_reg_22__retimed_I12746_QOUT;
reg x_reg_22__retimed_I12745_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12745_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845;
	end
assign N22149 = x_reg_22__retimed_I12745_QOUT;
reg x_reg_22__retimed_I12744_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12744_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061;
	end
assign N22147 = x_reg_22__retimed_I12744_QOUT;
reg x_reg_22__retimed_I12743_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12743_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627;
	end
assign N22145 = x_reg_22__retimed_I12743_QOUT;
reg x_reg_22__retimed_I12742_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12742_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967;
	end
assign N22141 = x_reg_22__retimed_I12742_QOUT;
reg x_reg_22__retimed_I12741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12741_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185;
	end
assign N22139 = x_reg_22__retimed_I12741_QOUT;
reg x_reg_22__retimed_I12740_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12740_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946;
	end
assign N22137 = x_reg_22__retimed_I12740_QOUT;
reg x_reg_22__retimed_I12739_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12739_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942;
	end
assign N22133 = x_reg_22__retimed_I12739_QOUT;
reg x_reg_22__retimed_I12738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12738_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681;
	end
assign N22131 = x_reg_22__retimed_I12738_QOUT;
reg x_reg_22__retimed_I12737_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12737_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919;
	end
assign N22129 = x_reg_22__retimed_I12737_QOUT;
reg x_reg_22__retimed_I12736_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12736_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532;
	end
assign N22125 = x_reg_22__retimed_I12736_QOUT;
reg x_reg_22__retimed_I12735_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12735_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942;
	end
assign N22123 = x_reg_22__retimed_I12735_QOUT;
reg x_reg_22__retimed_I12734_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12734_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777;
	end
assign N22121 = x_reg_22__retimed_I12734_QOUT;
reg x_reg_22__retimed_I12733_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12733_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688;
	end
assign N22117 = x_reg_22__retimed_I12733_QOUT;
reg x_reg_22__retimed_I12731_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12731_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918;
	end
assign N22113 = x_reg_22__retimed_I12731_QOUT;
reg x_reg_22__retimed_I12730_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12730_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289;
	end
assign N22109 = x_reg_22__retimed_I12730_QOUT;
reg x_reg_22__retimed_I12728_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12728_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587;
	end
assign N22105 = x_reg_22__retimed_I12728_QOUT;
reg x_reg_22__retimed_I12727_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12727_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571;
	end
assign N22101 = x_reg_22__retimed_I12727_QOUT;
reg x_reg_22__retimed_I12725_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12725_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813;
	end
assign N22097 = x_reg_22__retimed_I12725_QOUT;
reg x_reg_22__retimed_I12723_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12723_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028;
	end
assign N22091 = x_reg_22__retimed_I12723_QOUT;
reg x_reg_22__retimed_I12719_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12719_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909;
	end
assign N22082 = x_reg_22__retimed_I12719_QOUT;
reg x_reg_22__retimed_I12718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12718_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745;
	end
assign N22080 = x_reg_22__retimed_I12718_QOUT;
reg x_reg_22__retimed_I12715_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12715_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846;
	end
assign N22072 = x_reg_22__retimed_I12715_QOUT;
reg x_reg_22__retimed_I12713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12713_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049;
	end
assign N22066 = x_reg_22__retimed_I12713_QOUT;
reg x_reg_22__retimed_I12712_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12712_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296;
	end
assign N22064 = x_reg_22__retimed_I12712_QOUT;
reg x_reg_22__retimed_I12709_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12709_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169;
	end
assign N22056 = x_reg_22__retimed_I12709_QOUT;
reg x_reg_22__retimed_I12706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12706_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899;
	end
assign N22048 = x_reg_22__retimed_I12706_QOUT;
reg x_reg_22__retimed_I12703_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12703_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877;
	end
assign N22040 = x_reg_22__retimed_I12703_QOUT;
reg x_reg_22__retimed_I12701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12701_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[15];
	end
assign N22034 = x_reg_22__retimed_I12701_QOUT;
reg x_reg_22__retimed_I12690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12690_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[34];
	end
assign N22007 = x_reg_22__retimed_I12690_QOUT;
reg x_reg_22__retimed_I12689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12689_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[34];
	end
assign N22005 = x_reg_22__retimed_I12689_QOUT;
reg x_reg_22__retimed_I12688_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12688_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[16];
	end
assign N22003 = x_reg_22__retimed_I12688_QOUT;
reg x_reg_22__retimed_I12687_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12687_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[33];
	end
assign N21997 = x_reg_22__retimed_I12687_QOUT;
reg x_reg_22__retimed_I12685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12685_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[15];
	end
assign N21993 = x_reg_22__retimed_I12685_QOUT;
reg x_reg_22__retimed_I12682_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12682_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[12];
	end
assign N21983 = x_reg_22__retimed_I12682_QOUT;
reg x_reg_22__retimed_I12679_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12679_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[14];
	end
assign N21973 = x_reg_22__retimed_I12679_QOUT;
reg x_reg_22__retimed_I12676_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12676_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[11];
	end
assign N21963 = x_reg_22__retimed_I12676_QOUT;
reg x_reg_22__retimed_I12673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12673_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[13];
	end
assign N21953 = x_reg_22__retimed_I12673_QOUT;
reg x_reg_22__retimed_I12670_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12670_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[6];
	end
assign N21943 = x_reg_22__retimed_I12670_QOUT;
reg x_reg_22__retimed_I12667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12667_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[5];
	end
assign N21933 = x_reg_22__retimed_I12667_QOUT;
reg x_reg_22__retimed_I12664_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12664_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[8];
	end
assign N21923 = x_reg_22__retimed_I12664_QOUT;
reg x_reg_22__retimed_I12661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12661_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[10];
	end
assign N21913 = x_reg_22__retimed_I12661_QOUT;
reg x_reg_22__retimed_I12658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12658_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[7];
	end
assign N21903 = x_reg_22__retimed_I12658_QOUT;
reg x_reg_22__retimed_I12655_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12655_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[9];
	end
assign N21893 = x_reg_22__retimed_I12655_QOUT;
reg x_reg_22__retimed_I12652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12652_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[4];
	end
assign N21883 = x_reg_22__retimed_I12652_QOUT;
reg x_reg_22__retimed_I12649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12649_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[2];
	end
assign N21873 = x_reg_22__retimed_I12649_QOUT;
reg x_reg_22__retimed_I12646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12646_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[1];
	end
assign N21863 = x_reg_22__retimed_I12646_QOUT;
reg x_reg_22__retimed_I12643_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12643_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[3];
	end
assign N21853 = x_reg_22__retimed_I12643_QOUT;
reg x_reg_22__retimed_I12636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12636_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311;
	end
assign N21833 = x_reg_22__retimed_I12636_QOUT;
reg x_reg_22__retimed_I12635_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12635_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449;
	end
assign N21831 = x_reg_22__retimed_I12635_QOUT;
reg x_reg_22__retimed_I12632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12632_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171;
	end
assign N21818 = x_reg_22__retimed_I12632_QOUT;
reg x_reg_22__retimed_I12562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12562_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971;
	end
assign N21574 = x_reg_22__retimed_I12562_QOUT;
reg x_reg_22__retimed_I12560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12560_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108;
	end
assign N21570 = x_reg_22__retimed_I12560_QOUT;
reg x_reg_22__retimed_I12557_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12557_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327;
	end
assign N21559 = x_reg_22__retimed_I12557_QOUT;
reg x_reg_22__retimed_I12474_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12474_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162;
	end
assign N21310 = x_reg_22__retimed_I12474_QOUT;
reg x_reg_22__retimed_I12472_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12472_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300;
	end
assign N21306 = x_reg_22__retimed_I12472_QOUT;
reg x_reg_22__retimed_I12391_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12391_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439;
	end
assign N21064 = x_reg_22__retimed_I12391_QOUT;
reg x_reg_22__retimed_I12389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12389_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944;
	end
assign N21060 = x_reg_22__retimed_I12389_QOUT;
reg x_reg_22__retimed_I12340_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12340_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843;
	end
assign N20916 = x_reg_22__retimed_I12340_QOUT;
reg x_reg_22__retimed_I12338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12338_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977;
	end
assign N20912 = x_reg_22__retimed_I12338_QOUT;
reg x_reg_22__retimed_I12335_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12335_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194;
	end
assign N20903 = x_reg_22__retimed_I12335_QOUT;
reg x_reg_22__retimed_I12333_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12333_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334;
	end
assign N20899 = x_reg_22__retimed_I12333_QOUT;
reg x_reg_22__retimed_I12330_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12330_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920;
	end
assign N20890 = x_reg_22__retimed_I12330_QOUT;
reg x_reg_22__retimed_I12328_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12328_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054;
	end
assign N20886 = x_reg_22__retimed_I12328_QOUT;
reg x_reg_22__retimed_I12325_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12325_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275;
	end
assign N20876 = x_reg_22__retimed_I12325_QOUT;
reg x_reg_22__retimed_I12323_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12323_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414;
	end
assign N20872 = x_reg_22__retimed_I12323_QOUT;
reg x_reg_22__retimed_I12241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12241_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004;
	end
assign N20654 = x_reg_22__retimed_I12241_QOUT;
reg x_reg_22__retimed_I12232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12232_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086;
	end
assign N20632 = x_reg_22__retimed_I12232_QOUT;
reg x_reg_22__retimed_I12230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12230_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222;
	end
assign N20628 = x_reg_22__retimed_I12230_QOUT;
reg x_reg_22__retimed_I12229_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12229_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444;
	end
assign N20625 = x_reg_22__retimed_I12229_QOUT;
reg x_reg_22__retimed_I12227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12227_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950;
	end
assign N20621 = x_reg_22__retimed_I12227_QOUT;
reg x_reg_22__retimed_I12224_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12224_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168;
	end
assign N20613 = x_reg_22__retimed_I12224_QOUT;
reg x_reg_22__retimed_I12222_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12222_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306;
	end
assign N20609 = x_reg_22__retimed_I12222_QOUT;
reg x_reg_22__retimed_I12129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12129_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309;
	end
assign N20382 = x_reg_22__retimed_I12129_QOUT;
reg x_reg_22__retimed_I12124_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12124_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895;
	end
assign N20370 = x_reg_22__retimed_I12124_QOUT;
reg x_reg_22__retimed_I12118_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12118_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089;
	end
assign N20355 = x_reg_22__retimed_I12118_QOUT;
reg x_reg_22__retimed_I12103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12103_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872;
	end
assign N20295 = x_reg_22__retimed_I12103_QOUT;
reg x_reg_22__retimed_I12101_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12101_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829;
	end
assign N20290 = x_reg_22__retimed_I12101_QOUT;
reg x_reg_22__retimed_I12099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12099_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040;
	end
assign N20285 = x_reg_22__retimed_I12099_QOUT;
reg x_reg_22__retimed_I12097_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12097_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063;
	end
assign N20280 = x_reg_22__retimed_I12097_QOUT;
reg x_reg_22__retimed_I12095_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12095_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259;
	end
assign N20275 = x_reg_22__retimed_I12095_QOUT;
reg x_reg_22__retimed_I12093_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12093_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285;
	end
assign N20270 = x_reg_22__retimed_I12093_QOUT;
reg x_reg_22__retimed_I12091_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12091_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234;
	end
assign N20265 = x_reg_22__retimed_I12091_QOUT;
reg x_reg_22__retimed_I12089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12089_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852;
	end
assign N20260 = x_reg_22__retimed_I12089_QOUT;
reg x_reg_7__retimed_I11924_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I11924_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367;
	end
assign N19755 = x_reg_7__retimed_I11924_QOUT;
reg x_reg_7__retimed_I11922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I11922_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869;
	end
assign N19751 = x_reg_7__retimed_I11922_QOUT;
reg x_reg_7__retimed_I11834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I11834_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317;
	end
assign N19431 = x_reg_7__retimed_I11834_QOUT;
reg x_reg_7__retimed_I11739_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I11739_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22];
	end
assign N19158 = x_reg_7__retimed_I11739_QOUT;
reg x_reg_26__retimed_I11459_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__retimed_I11459_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594;
	end
assign N18406 = x_reg_26__retimed_I11459_QOUT;
reg x_reg_26__retimed_I11457_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__retimed_I11457_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897;
	end
assign N18402 = x_reg_26__retimed_I11457_QOUT;
reg x_reg_22__retimed_I11390_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I11390_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82;
	end
assign N18245 = x_reg_22__retimed_I11390_QOUT;
reg x_reg_22__retimed_I11388_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I11388_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741;
	end
assign N18241 = x_reg_22__retimed_I11388_QOUT;
assign N22961 = !N18241;
assign N22966 = !N22961;
assign N22965 = !N22961;
assign N22964 = !N22961;
assign N22963 = !N22961;
assign N22962 = !N22961;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161 = !(a_exp[7] & a_exp[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854 = !((a_exp[6] & a_exp[5]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13163);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13161 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18854);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18861;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201 = !(((a_man[0] | a_man[1]) | a_man[2]) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13197);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212 = !(a_man[4] | a_man[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13184 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13203) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13192) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13212);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24 = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13201) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13195) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13206) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13216);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__19 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__24;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110 = ((a_exp[7] | a_exp[6]) | a_exp[0]) | a_exp[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114 = ((a_exp[4] | a_exp[2]) | a_exp[3]) | a_exp[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13110 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13114);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141 = !(((a_exp[1] & a_exp[2]) | a_exp[3]) | a_exp[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138 = !((a_exp[6] & a_exp[5]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13141));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21 = !(a_exp[7] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13138));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385 = !a_exp[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364 = !a_exp[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373 = !(a_exp[2] & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371 = a_exp[4] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379 = a_exp[5] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376 = !(a_exp[6] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376 ^ a_exp[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5379 ^ a_exp[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5376 | (!a_exp[7]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18845 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__17 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__21) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__46;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N741;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13910;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N594));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612 = !a_man[21];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270} = {1'B0, a_man[22]} + {1'B0, a_man[20]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957} = {1'B0, a_man[21]} + {1'B0, a_man[19]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042} = {1'B0, a_man[22]} + {1'B0, a_man[19]} + {1'B0, a_man[17]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361} = {1'B0, a_man[20]} + {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4204};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391} = {1'B0, a_man[18]} + {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4545} + {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4042};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612 | a_man[19];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185} = {1'B0, a_man[17]} + {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4506};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198 = !a_man[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198 | a_man[20];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4170} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4229} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4391};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198) ^ a_man[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291 = !a_man[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291 | a_man[18];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081} = {1'B0, a_man[16]} + {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4130};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4571} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4185};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612) ^ a_man[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975 = !a_man[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975 | a_man[17];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976} = {1'B0, a_man[15]} + {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4466};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4193} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4348} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4081};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291) ^ a_man[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385 = !a_man[18];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385} + {1'B0, a_man[13]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594} = {1'B0, a_man[14]} + {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4404};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4533} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3970} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3976};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975) ^ a_man[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069 = !a_man[17];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183} = {1'B0, a_man[12]} + {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588} = {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4336} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4029};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4158} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4311} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4594};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471 = !a_man[16];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4588} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3960} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4183};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4092} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4246} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4488};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565 = !a_man[14];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420} = {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162 = !a_man[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359} = {1'B0, a_man[22]} + {1'B0, a_man[13]} + {1'B0, a_man[10]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4232} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4577} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4359};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006} = {1'B0, a_man[11]} + {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4300};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4455} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4395} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4126};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4521} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4428} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4617};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377} = {1'B0, a_man[12]} + {1'B0, a_man[9]} + {1'B0, a_man[7]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161} = {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625} = {1'B0, a_man[8]} + {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4314};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4510} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4420} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4377};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4324} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4173};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4207} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4365} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4006};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253 = !a_man[13];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288} = {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031} = {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135} = {1'B0, a_man[7]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4186};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4383} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4609} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4625};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4444} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4043} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4351};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4078} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4147} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4241};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939 = !a_man[12];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630} = {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368} = {1'B0, a_man[6]} + {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4058};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4252} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4470} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4135};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4288} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4640} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4221};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4264} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4018} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4260};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339 = !a_man[11];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613} = {1'B0, a_man[5]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4630};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4120} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4338} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4368};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4161} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4500} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4093};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4137} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4197} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4495};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032 = !a_man[10];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4210} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4236} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4613};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4031} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4369} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3963};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4002} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4067} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4016};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474} = {1'B0, a_man[6]} + {1'B0, a_man[3]} + {1'B0, a_man[1]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121 = !a_man[8];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601} = {1'B0, a_man[22]} + {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4266} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4023} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4237};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432 = !a_man[9];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432} + {1'B0, a_man[4]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4200} + {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4123};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3987} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4082} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4549};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4591} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3936} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4249};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525 = !a_man[7];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4046} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4386} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4601};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473} = {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621} = {1'B0, a_man[5]} + {1'B0, a_man[2]} + {1'B0, a_man[0]};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4138} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4641} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4474};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4107} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4653};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4524} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4457} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4485};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097 = !a_man[6];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940} = {1'B0, a_man[13]} + {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4187} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4096} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4012};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4473} + {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4621};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3977} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4421};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4486} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4397} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4004};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631 = !a_man[5];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247} = {1'B0, a_man[1]} + {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4372};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4566} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4541} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4070};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4614} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3952} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4355};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175} = {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511} = {1'B0, a_man[3]} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4655};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4124} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4033} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4247};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4306} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4211} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4511};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4458} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3940} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3965};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4317} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4409} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4493};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445 = !a_man[3];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4049} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3955} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4175};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304 = !a_man[4];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086} = {1'B0, a_man[2]} + {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4056};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4400} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4489} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4238};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4255} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4597} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4132};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410} = {1'B0, a_man[1]} + {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4227};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4423} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4331} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4086};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4527} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4151} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4394};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398 = !a_man[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505 = a_man[15] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4505};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3980} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4618} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4410};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4166} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4073} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3953};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4320} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4516} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4543};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4179} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4268} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3937};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333 = (!a_man[15]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4214} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4284} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4333};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434 = !a_man[1];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4215};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4258} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4346} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4100};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4110} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4449} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4293};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244} = {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4198};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4156} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4403} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4574};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4129} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4191};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4009} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4388} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4550};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966 = !a_man[0];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353} = {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4116} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4335} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4244};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4064} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3993};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4037} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3944} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4101};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592} = {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4427} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4519} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4353};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4586} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4182};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3969} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4636} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4454};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4291};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109} = {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4624} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3984} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4592};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4052} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4364};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4090} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4556} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4000};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3975};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343} = {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4385} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4076} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4172} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4109};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4230} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4546};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4271} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4027} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4235};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4638);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104 = a_man[9] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948 = (!a_man[9]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3948};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4104} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4649};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4206} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4453} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4472};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4069};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4041} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4507} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4343};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4393} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4014} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3988};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4001);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4471} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4536} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4219} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4360};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4608} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4573} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4225};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4480;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4145;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498 = a_man[5] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4498};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4162};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4066} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4160};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4639} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4382} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4478};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4287} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4442} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4242};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4565} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3999} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4560} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4604};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626} = {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4253} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337 = (!a_man[5]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4337} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4184} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3995};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136} = {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4339};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015} = {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3962} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4015};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4429} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4626};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4456} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4250};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4208} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4136};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4121} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4396} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4367};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4525} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4097};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4484} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4234};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4325};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966} + {1'B0, a_man[6]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4445;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978 = !(a_man[1] | a_man[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4398;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3966 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4290);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4088 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4402) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4243);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3978) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4201)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4047);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4434 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4199);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4513 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4352);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4554 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4154;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4308 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3992) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4329) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4514);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4634) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4595)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3950) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4021));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4174 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4652);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4222 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4213) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4062);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4530) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4580)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4080) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4548));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3985 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4148);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4301 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4628);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3968 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4282;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4437 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4127) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4118) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4563);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4576) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4508);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4055 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4366);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4522 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4117);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4344) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4190);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4274 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4590);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4030 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4248);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4503 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4256) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4098);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4418) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4481)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4323);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4283 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4600;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4406 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4467 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3972);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4413 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4007;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4165 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4567) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4347) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3961);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4134 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4194);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4350 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4322);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4318 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4071) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4643);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4460) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4529)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4373);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18828) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3935)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18830) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18832));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4298 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3958);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4559 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4312) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4114 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4494)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4128) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4602)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4439);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4658 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4309);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4468 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4220) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4463 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4438)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4603 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4414);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4569 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4141)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4504)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4345);
assign N22968 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4025;
assign N22971 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4178 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422);
assign N22969 = !(N22968 & N22971);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059 = !N22969;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4295 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4584);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4024 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4552)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3989 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4280);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4433 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4005)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4415)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4257);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4163 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4292);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4447 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4177)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4326 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4149);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4302 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4276)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4319)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4167);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4085) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4526)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4371);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4430 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4407);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4562 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4538)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3974 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3949);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4105 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4482)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4226)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4072);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4651 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4627);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4053 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4115)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4496);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4557 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3934)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4142)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3979);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3990 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4341);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3996 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4218);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4378 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4605)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4039 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4262);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4417 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4647)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4048)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4619);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4297 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4075);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4451 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4622)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4361 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4051);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464) | (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3957 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4518)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3954)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4515);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4632) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4459);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4435)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4279);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4112 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4270);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4612 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4425) & (!(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376)));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4499);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169 = (!a_man[22]) ^ a_man[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4139;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4635;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3946)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4102);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4261) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4376;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3938 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4169) & (a_man[22] | a_man[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1] = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5364;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N37297;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4356;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4305;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4150;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4223)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4387);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4202;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4119) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4275);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4540;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4089;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4217)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4380);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4532) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4555;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4606 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4063;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4155;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3994;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4431) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4440)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4607);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4038) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4464;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[1] ^ a_exp[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5373 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5385;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5371) ^ a_exp[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5372 ^ a_exp[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N650) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N651));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N652 & a_exp[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N646) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N647));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N648) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N649));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5578 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N706) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5585) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5491));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4441 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4245;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4448;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4501;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4294;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4629) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4057);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4181;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3998)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4157);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4310) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4657;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5612) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5464 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5606 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N704;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4209 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4334;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4216;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4272;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4497)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3933);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4091) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4028;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5519) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5434));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5409 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5513 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N702) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N644) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N645));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5443) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4285 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4426;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N641));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N642) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N643));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5512 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5416) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5540));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5465 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N701) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5565) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5473));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5482));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5455 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5558 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N703;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5577));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5598 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5436 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N705;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6280;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6209 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6355);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6125 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5921 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178 = 1'B0 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6470 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6057 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6478 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6254);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[27] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5965 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6172 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[27]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6003 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5890 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6332 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6103 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6251 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[26] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6519 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6022 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[26]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6066 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6446 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6175 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5952);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5940 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5936 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[25] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6369 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6564 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[25]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4399) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4239);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4542)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4389);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4363);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4587 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4113;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3986) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4520;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5594) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5511));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5568) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5580 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N699) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4316;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4452);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3959 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4205;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N638));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N639) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N640));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5462));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5521) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5485 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N698) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5425) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5546));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5557));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5531) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5417 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N700 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8912;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42] = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9401 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6042);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N763;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8700) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6299 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6024 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6507 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6493 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6488 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[24] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6217 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6412 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[24]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6144 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6567 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6189 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6341 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[23] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6067 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6265 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[41] = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[42];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4131) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4623;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N637));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5499) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5415));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5474) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5560 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5494 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5604) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5608));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N697) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4596;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4645)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4476);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4547);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4054 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4299;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N636));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5450) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5584));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5427) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5444 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5467 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5616 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5509) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5515));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N696) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8946;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9435 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8724) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6431 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6491 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5970 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6566 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N762;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8752) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[41], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[40]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9092};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[41]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[23]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[41]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6415 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6494 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6134 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6580 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6185 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[22] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5897 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6110 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6285 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6342 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6523 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6414 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N761;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8811) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9628;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8779) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4083) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3983;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N635));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5405) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5538));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5597) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5613 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5587 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5523 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5414) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5419));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N695) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4065;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4648);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4146 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4392;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5574) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5549) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5566 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5493 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5428 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5537) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5542));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N694) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8982;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6239 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6178 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6131 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6188 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6376 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6267 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N760;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8871) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9128} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10066};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[40], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[39]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9236} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8732} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9847};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[22]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[40]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[40]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144 = N22678 & N22680;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6088 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6268 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6427 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6036 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[21] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6453 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5948 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9468 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8748) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3971) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4077;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N633));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5442));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5503) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5520 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5446 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5550 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5440) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5447));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N693) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4008;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4490;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4330;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4095)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4254);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4568;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4582) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4022);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4013;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4650)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4079);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4231) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4479;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N632));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5479) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5611));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5453) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5472 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5615 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5456 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5569));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N692) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9013;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8842) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9555} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8766};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8902) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8807) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9166} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10100} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9163};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6090 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6028 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6168 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5971 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6038 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6223 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6112 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N759;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8935) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9707} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8986} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8924};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[39], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[38]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9302} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9467} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10055};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[39]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[39]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6113 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6440 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6282 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6577 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[20] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6308 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6502 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9497 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8776) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4176 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4171;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N631));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5431) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5564));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5406) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5461));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5424 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5470) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5476));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N691) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4411;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4103;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4419)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4579);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4017) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4575;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N630));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5601) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5518));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5576) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5413));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5595 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5591) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5599));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N690) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9050;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6212 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6207 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5922 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6571 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6525 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6579 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5950 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N758;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6061 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6475 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6417 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6560 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6074 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6426 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5903 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6505 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N757;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9057) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9595} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8940};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8997) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9321} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8699} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8648};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8869) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6329 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6270 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6279 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6456 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6360 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N756;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9122) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8840) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9200} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8609} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9228};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8797} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9742} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8624};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9024) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8932) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9528 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8805) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4534 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4263;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N629));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5553) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5471));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5530) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5583));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5547 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5497) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5505));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N689) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4099)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3945);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4195);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4509 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3947;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N628));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5507) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5422));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5481) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5535));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5402) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5408));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N688) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9086;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9087) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9630} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8974};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10135} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9358} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10210};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10088} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9045};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9438} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10114} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10178};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[38], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[37]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8774} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9691} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9529};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[38]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[38]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6474 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5951 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6343 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6424 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[19] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6153 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6356 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8899) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6444 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6173 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6116 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6458 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6124 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6312 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6202 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N755;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9188) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8995) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9920} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8834} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9781};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9247} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9940} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9724};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9218) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5892 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6304 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6023 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5955 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6182 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6314 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5964 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6159 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6049 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N754;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6565 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6509 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6160 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6518 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6000 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5882 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N753;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9323) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8929) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9158} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9956} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8866};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9562 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8836) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3951) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4349;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N627));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5459) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5403) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5592));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5433) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5487));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5452 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5525) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N687) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4059;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4286);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4611 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4040;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5411) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5571) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5545));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5602) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5441));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5404 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5430) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5435));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N686) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9124;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9118) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9668} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9005};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9256) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8867) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9242} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9546} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9294};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8758} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9510} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9974};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8961) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9153) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9055) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8638} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10173} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9392};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8656} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10123} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9854};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8870} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9149} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9637};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10002} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9019} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8751};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9109} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9818} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9883};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7328} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7459} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7293};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7375} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7822} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7709};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7344} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7316} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7896};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7887} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7473} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7682};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7753} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7616} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7751};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7787} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7543} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7608};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7322} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7300} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7455};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7837} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7734} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7592};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7872} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7471} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7330};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7926} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7909} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7687};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7665} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7817} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7878};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7395} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7676} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7308};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7731} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7697} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7835};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7379} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7527} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7538};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7754} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7535} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7814};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7452} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7556} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7411};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7765} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7626} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7745};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7599} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7761} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7337};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7893} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7903} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7314};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7465} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7613} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7924};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7545} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7702} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7841};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7838} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7620} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7476};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7388} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7925} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7775};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7680} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7911} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7483};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7325} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7639} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7394};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7336} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7341} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7828};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7780} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7417} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7560};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7927} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7699} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7557};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7900} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7499} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7640};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7694} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7354} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7826};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7628} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7365} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7865};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7759} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7342} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7730};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7503} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7643} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7931};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7356} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7777} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7641};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7333} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7859} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7355};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4379) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4443;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N625));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5581) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5486));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5526) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5498));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5554) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5610));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5552) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5556));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N685) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7918} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7706} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7407};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7720} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7549} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7480};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7843} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7667} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7301};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7707} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7451} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7358};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7586} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7726} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7359};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7440} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7861} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7723};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7414} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7581} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7722};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4535;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4192;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4036;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4422 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4446) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4615);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4381;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4045) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4384)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4537);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N3973) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N4133;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438 = !((a_exp[0] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N623) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N624));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5534) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5438));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5478) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5500) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5449));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5510) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5562));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5528 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5423);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5458) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5463));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N684 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5817;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7437} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7915} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7565};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7421} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7813} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7725};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7830} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7746} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7380};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7526} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7806} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7444};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7524} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7297} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7804};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7500} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7296} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7438};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7908) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7770;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7785} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7534};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7520} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7562} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7494};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7552} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7692} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7635};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7800} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7625};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7920} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7611} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7891};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7609} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7378} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7888};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7582} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7661} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7801};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7790);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7882} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7507};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7339} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7522} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7346};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7442} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7349} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7405} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7492} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7769};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7688} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7464} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7323};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7663} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7377} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7523};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7576} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7604} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7885};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7795} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7852} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7574};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7712} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7705};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7899} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7805} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7431};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7766} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7402} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7550};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7744} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7742} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7886};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7869} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7619} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7525};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7419} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7606};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7517} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7290} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7657};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7849} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7633} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7488};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7827} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7463} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7607};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7369);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7684} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7320};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7889} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7880} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7372};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7426} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7319} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7332};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7286} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7572} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7713};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7825} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7916} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7321};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7306} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7791} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7782};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7698} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7610} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7739};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7370} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7792} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7655};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7547} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7347} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7686};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7876);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7505} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7513} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7398};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7413} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7324};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7736} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7457} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7877};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7428} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7914} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7400};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7399} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7763} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7875};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7867} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7776};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7819} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7540} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7597};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7630} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7514} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7764};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7588} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7596};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7690} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7906} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7679};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7312} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7345} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7486};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7304} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7860} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7768};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7595);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7456);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7845} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7311};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7484} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7404} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7623};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7757} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7424} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7569};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7710} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7392} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7847};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7310);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7670} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7568};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7788} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7479} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7938};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7818);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7935} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7391};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7490} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7509} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7650};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7383} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7851} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7366};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7678);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7749} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7648};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7539);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7364} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7469};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7669) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7482)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7386));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7532 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7672);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7600 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7303) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7808);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7587) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7430)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7811) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7307));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7448 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7591);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7829 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7866) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7504) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7585)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7729) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7870));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7363 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7508);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7905 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7781) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7645);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7647 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7786);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7936 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7933 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7704) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7563);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7571) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7632)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7487);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7567 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7708);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7844 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7343);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7485 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7629);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7762 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7912);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7397 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7546);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7685 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7824);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7318 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7462);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7603 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7741);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7883 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7374);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7519 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7659);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7797 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7292);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7434 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7577);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7854 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7718);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7495 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7351);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7637 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7772);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7408 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7922);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7554 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7695);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7327 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7832);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7614 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7468);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7601 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7748);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7302) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7807;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7689) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7425) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7939;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7812) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7674;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7427 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7940));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[32] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7409 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7443;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7580;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7660;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7376) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7884;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7521 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7294) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7799;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7436 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7858) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7719;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7668) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7528;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7403) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7917;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7789) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7652;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7533) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7387;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7566 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7420));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7773 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7666;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[32]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10143;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9397;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[37], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[36]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9140} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9208} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10121};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[37]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[37]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6187 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6286 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6326 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6506 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6264 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5967 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6277 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[18] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5995 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6199 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[19] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9286) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8894) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9276} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9588} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9362};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9020) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8991) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9185) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9084) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8668} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10206} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9432};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9813} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9091} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8875};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9596 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[3]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8864) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9150) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9702} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9040};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5939 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5986 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6413 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6363 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6274 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6002 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6368 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6550 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6438 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N752;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9388) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9254) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9353) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8958) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9195} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9988} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8901};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8789} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9455} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10192};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10094} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9119} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9644};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9763} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8579} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9283};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6266 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6205 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6120 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6552 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6216 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6398 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N751;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9457) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9051) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[1] & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923 | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8892) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8956) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9694} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9350};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8927) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9315} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9841} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7288};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9851} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10128} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10018};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9223} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8731} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10216};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8678} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9889} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8907};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8782} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9539} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10038};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9912} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8674} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8934};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6405);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6020 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5975);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[18] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9502} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9790} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8855};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[36], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[35]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8839} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9620} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8897};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[18]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[36]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[36]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12300;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7467;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7636;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7796;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7317;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7396 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7910;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7823 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7881) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7740;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7658 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7717) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7575;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7493 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7553) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7406;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7326 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7381) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7892;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7767) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7634;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7511) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7368;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7897) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7752;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7934 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7784));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7496 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7890;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7831;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7350;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7518;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7544 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7602) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7460;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7373 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7432) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7291;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7853 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7921) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7771;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7693 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7747) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7612;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7489) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7348;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7874) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7733;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7617) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7472;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7646 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7506));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7855 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7466;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9524 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5945 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6495 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[17] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6536 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6425 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9115) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6111 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6054 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5958 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6065 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6248 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6137 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N750;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9520) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9419) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9772} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9470} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8826};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9215) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9319) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9018) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9621} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8692} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10237};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9805} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8825} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9063};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9182) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9736) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9660;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6472 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5949 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5885 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6513 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6377 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6098 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5896 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6096 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5979 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N749;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9590) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9459} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9077} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9386};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9284) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9384) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8988) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9231} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10027} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8937};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9654} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9623} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8667};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9832} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9587} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8849};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9979} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9255} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9002};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9487) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9081) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9349) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9251) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9269} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9661} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8723};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9884} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10164} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8694};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9425} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9391} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10163};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9615} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8640} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8661};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10008} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9771} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9027};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9415} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9674} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10158};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6316 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6345 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6053);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[16] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6385 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6123 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8601} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9056} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9066};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9407} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9837} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9699};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[35], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[34]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10233} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8810};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6171 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6361 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6520 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6122 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[17] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6547 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6046 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12171} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[17]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[35]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[35]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838 = !(N21831 & N21833);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5957 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6479 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6017 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6203 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6354 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6371 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5961 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[16] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6395 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5879 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[31]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10180;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[30]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8922) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6161 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6192 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6293 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5884 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6358 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[15] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6232 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5963 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9552) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9048) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6503 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6443 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6225 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5934 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6452 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5933 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N748;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9656) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8603} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9806} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9000};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9431} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9230} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9987};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9194} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10137} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9955};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6357 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6296 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6529 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6210 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6075 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6307 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6481 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6382 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N747;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9716) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9112) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9518) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9915} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8662} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10197};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9316) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9416) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8595));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9016) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9267} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10058} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8970};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10208} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9241} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10026};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9454) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9146) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9212) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9775) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9618) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9305} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9114} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9422};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9504} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8857} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9469};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10172} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9203} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9008};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6200 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6142 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6058);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5907 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6154 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6033 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6152 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6339 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6229 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N746;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9782) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9282) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9179) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8753} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9980} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9541};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9381) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8754;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9693} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10145};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9907));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9079) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9684) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8632} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9842} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9031};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9727} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9503} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10236};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9039} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9997} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9814};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9780} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9964} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8796};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9165} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8973} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9928};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9357} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9385} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10099};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7624) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7481;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7313 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7793;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7287 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7458) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7537);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7447 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7305));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7352) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7491;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7338) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7842;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7681 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7515;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7656 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7820) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7902);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7810 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7671));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7857) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7715;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7907) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7758;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7598 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7429;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7737) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7816);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7728 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7590));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7498) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7919;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9325 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9797} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8788} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8706} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10047} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9186};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7371;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7703;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7541) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7393;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7879 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7850) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7714;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7594) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7454;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7331) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7836;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7362 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7868));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7578 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7691;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9424 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10061} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9824} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9311};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[34], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[33]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9996} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10150} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8726};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897} = {1'B0, N22003} + {1'B0, N22005} + {1'B0, N22007};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032 & N21818);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9627 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8984) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9043) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[29]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9248;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[28]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8832) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8845, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10185} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9047} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9238} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9447};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[33], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[32]} = {1'B0, N22145} + {1'B0, N22147} + {1'B0, N22149};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6056 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6025 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6562 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6050 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6521 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6351 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6007 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6219 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6515 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[15] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6435 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251} = {1'B0, N21993} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[33]} + {1'B0, N21997};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6517 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6410 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5883 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6102 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6218 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6068 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6366 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[14] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6093 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6288 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6006 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6211 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6442 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6201 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[14] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6085 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6516 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8889) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9946, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9578} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9292} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8817} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8698};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9108) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6253 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6335 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6582 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6295 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6048 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[13] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5917 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6367 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9078} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9850} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8865};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9747) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9144) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9947} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8686} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10230};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8602} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9343} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9113};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9451) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9249) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8784;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9151} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9306} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10205};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9484) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9652) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9347) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5966 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6047 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5984 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6574 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5994 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6181 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6082 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N745;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9843) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10090} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9460} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9613};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8891} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9766} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9540};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9277} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10034} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9631};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9015} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8833} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9788};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6141 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6076 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5880 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6538 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6421 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6546 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6031 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5913 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N744;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9905) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9313) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9811) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8785} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10016};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9527);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9413) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9226} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9728};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9714) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9616) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9515) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9877} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9067} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8928};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9800} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8820} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9581};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9885} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9314} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8900};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8672} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9049} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9398};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9594} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8644} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8803};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8981} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9557} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9751};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7299 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7756) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7622);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7531 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7385));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7721) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7289;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7932 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7478) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7895 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7750));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7579) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7516;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9220 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9744} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8949} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10130} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8590} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9129};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8953) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[27]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10039;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[26]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8741) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9176) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9919} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9856} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10031} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10203};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8967, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8629} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9548} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8863} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8608};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[32], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[31]} = {1'B0, N22137} + {1'B0, N22139} + {1'B0, N22141};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976} = {1'B0, N21973} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[32]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[32]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839 = N20872 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6224 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6302 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6250 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6428 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6387 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6167 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6337 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6140 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5881 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[12] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6467 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6215 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8799) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9523} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8765} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9475};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6100 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6283 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6400 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6179 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6359 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5983 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6437 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[11] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6324 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6063 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9379} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9152} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9914};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9875) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9378) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9778) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10124} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9655} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8717};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9617} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9418} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10160};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9278) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9835;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10193} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9190} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8772) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9136));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9210) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9682) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9482) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6261 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5878 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6436 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6388 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6578 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6301 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6094 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6272 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6394 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6464 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N743;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9342} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9496} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8850};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9582} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9064} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8852};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8631} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9352} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8936};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10063} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9667} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9085};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9933) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5941 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6289 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6235 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6146 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6119 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6420 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6320 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N742;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10028) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10190} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9262} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8649};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9583) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9344) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9448) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9839) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9764} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8818} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10050};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8597} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10075} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9873};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9189} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8663} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9950};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9701} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10096} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8728};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8701} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9857} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9440};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9819} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10147} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8841};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7644 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7840) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7701);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7615 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7470));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7435) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7738;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7627 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7559) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7416);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7329 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7833));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7295) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7315;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9121 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9363} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9564} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8769} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8613} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8770};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9012) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9245) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8587} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9666} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9715} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9849};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9320, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8942} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9157} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9896} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8911};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[31], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[30]} = {1'B0, N22153} + {1'B0, N22155} + {1'B0, N22157};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6510 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6262 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6439 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6466 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6101 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5899 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6213 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[13] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5927 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6135 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335} = {1'B0, N21953} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[31]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[31]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[25]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9090;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[24]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8664) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8859) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9075) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10073} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9083} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8906} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9274};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9309) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6149 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5988 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5935 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6128 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6537 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6290 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[10] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6166 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5895 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8920) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9749} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10108} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8727};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9098} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9466} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9329} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9525};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9681, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9289} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8740} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9519} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9491};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[30], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[29]} = {1'B0, N22129} + {1'B0, N22131} + {1'B0, N22133};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6037 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6108 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6292 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5937 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6454 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[12] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6480 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5976 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055} = {1'B0, N21983} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[30]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[30]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9139) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8712) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6009 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6404 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6221 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6486 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5968 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6259 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6183 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6386 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[9] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6013 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6451 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9745) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9648) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9545) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9910} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9104} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8962};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8885} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8713} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10194};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9710) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9511) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9994) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9380} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9533} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8881};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10112);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9290);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10168) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10084) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9036} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8714} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9833};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9902) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9410) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9808) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10161} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9686} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8744};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10111} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9135} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9906};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9225} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9657} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9983};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9389} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8969} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10131};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9717} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9493} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10225};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9579) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9680) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10113) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8886} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8915} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9870};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9941} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8998} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9971};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9752} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8957} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8771};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9330) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10023) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10054) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8689));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9753);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9683} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10224} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9297};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9612) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9872) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9366));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9478) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9776) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9801} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10083} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9141};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8626} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9175} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9937};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8921} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9689} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9264};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8688} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9003} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9426};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9735} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9159} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8760};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9123} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9479} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9891};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7605 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7929) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7779);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7696 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7555));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7798) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7542;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7410 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7923));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7502 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7760;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9021 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21];
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10181} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8872} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8979} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9173} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9600};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8592, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8580} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8896} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8619};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869} = {1'B0, N22233} + {1'B0, N22235} + {1'B0, N22237};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[29], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[28]} = {1'B0, N22105} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10223} + {1'B0, N22109};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5974 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5905 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5947 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6447 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5900 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6012 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6489 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6309 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5893 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[11] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6333 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6530 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413} = {1'B0, N21963} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[29]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[29]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9445) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8767) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9720} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9888} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8722} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9935};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9275) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5888 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6237 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6184 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6373 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6541 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6086 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6531 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[7] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6407 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6151 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5924 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6391 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6071 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6340 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6522 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5990 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6408 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6016 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6234 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5977 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[8] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6558 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6306 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9836) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9929) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9645) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9721} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8778} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8657};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9741) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9542) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10025) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9417} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9572} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8919};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8992} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9759} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8806};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9526} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9722} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8594};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10021} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8719} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9034};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9774} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10166} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8791};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7774 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7638));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7863 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7340;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18] & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9923} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9513} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10212} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9199} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8908};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8828) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9639} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9882} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9509};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9041) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9960} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9209} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9697};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[23]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9895;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[22]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8585) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8983) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9207) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10060} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9706} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10235};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8745} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8651} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9370} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8954};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10049, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9688} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10082} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9903} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9103};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9375) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9296, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8918} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9074} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9336} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9133};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[28], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[27]} = {1'B0, N22064} + {1'B0, N22066} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9869};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6077 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6117 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6499 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5980 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6186 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6155 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6449 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[10] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6176 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6379 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137} = {1'B0, N21913} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[28]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[28]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9508) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8637) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[21]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8947;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[20]) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10157) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9106) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8685) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9312} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8763} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8941};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10117, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9322} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10057} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8675};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9341) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8884) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9576) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9120} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9500} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9690};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9143, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8777} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9969} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9409} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8989};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495} = {1'B0, N22249} + {1'B0, N22251} + {1'B0, N22253};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[27], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[26]} = {1'B0, N22113} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9879} + {1'B0, N22117};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6568 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6145 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5898 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6352 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6534 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6310 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5997 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6305 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[9] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6026 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6226 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864} = {1'B0, N21893} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[27]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[27]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9900) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9990) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9804) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9333} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10118} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9181};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8742} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9131};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8985);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10080) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9898} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9611} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8591};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9794} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8814} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9602};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9566} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8622} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8780};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9299} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8746} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10053};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7497 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7353));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7584) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7564;
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9462} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9809};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6190 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6581 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6576 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6069 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6240 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6043 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6511 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6532 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6469 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[5] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6106 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6206 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6035 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6220 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5918 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6380 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[6] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6256 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5993 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9197} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9551} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9427};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10170} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8943} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8581};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10215) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9174) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8739) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8933} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10101} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8606};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9250} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9676} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8708};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9406) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8951) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9643) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8757} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9111} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9304};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8813} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9449} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10004} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9022};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9909, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9532} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10152} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9757} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9180};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[26], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[25]} = {1'B0, N22080} + {1'B0, N22082} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9495};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6004 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6294 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6197 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6383 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6278 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6548 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6150 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[8] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6569 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6078 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215} = {1'B0, N21923} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[26]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[26]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8646));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9610) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9708) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9364);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9874) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10146) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10228));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10052) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9904} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9221} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8955};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9977} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9028} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8658};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8653} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9575} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9373};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9535} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9337} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10085};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9963} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9499} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9072};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5928 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6553 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5996 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6423 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5901 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5915 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6260 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6325 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6079 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[4] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5944 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6393 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10201} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8829} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8691};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10062) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9243) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9556} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9958} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8600};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8795) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8607) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9476) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9743} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9921} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8750};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9827} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9709} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9285} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8733};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9010) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10093} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8610} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8926};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8846} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9486} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10040} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9058};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9942, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9571} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10186} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9792} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9217};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[25], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[24]} = {1'B0, N22121} + {1'B0, N22123} + {1'B0, N22125};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5942 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6045 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6230 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5908 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5998 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6346 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6315 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6396 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5991 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[7] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5909 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943} = {1'B0, N21903} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[25]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[25]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8856) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8660) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9538) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9356} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9547} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10087};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9959) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9773) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9868) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9609} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9756} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8812};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9383} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9411} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10155};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8627} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10119} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9145};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8598} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9201} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9107};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5891 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6015 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6276 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6455 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5923);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6228 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6559 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5910 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[3] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6496 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6243 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10231} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9845} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9659};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8781));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10125) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9307) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9164} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9234} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9913};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10217, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9862} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8977} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9746} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9324};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9071) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9769) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9733} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9591} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8596};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9257, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8877} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8768} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10068} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9093};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608} = {1'B0, N22217} + {1'B0, N22219} + {1'B0, N22221};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[24], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[23]} = {1'B0, N22097} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9976} + {1'B0, N22101};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5877 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6127 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6401 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5876 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6083 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6460 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6193 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6246 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6543 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[6] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6269 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6462 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299} = {1'B0, N21943} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[24]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[24]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8917) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8711) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9607) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9156} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9726};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10110) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10022) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10104} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8620} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9371};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9967));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9677) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9738) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9927) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9834) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10153} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10009} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9216};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8680} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9192} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9952};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10126} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9183} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9944};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9346} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10174} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9911};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6051 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6389 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6104 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6121 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6311 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6139 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6055 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6081 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6227 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6463 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[2] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6348 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6092 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9308} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9880} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8887};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10120));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10188) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9372) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8798} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9270} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9537};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9521, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9130} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9991} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8641};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9134) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9830) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9348} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8860} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9908};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8588, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9899} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9784} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9360} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10103};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646} = {1'B0, N22209} + {1'B0, N22211} + {1'B0, N22213};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[23], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[22]} = {1'B0, N22072} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10011} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9608};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6459 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6191 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6434 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6303 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6328 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6095 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6392 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[5] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6114 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019} = {1'B0, N21933} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[23]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[23]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8980) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8764) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9675) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8639} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8790} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9340};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9760));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8582) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9802) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10076) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9986) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8990} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9647} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9793};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9598);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9399);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9718) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10175) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10077));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8617} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9359} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9936};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8793} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9553} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8822};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9978} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8999} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8972};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9155} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9430} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8965};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10141) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9206);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10048) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8642} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8650} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9408};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9897) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8847} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9901} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10132};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9585} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8611} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8635};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9768} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8787} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9739};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9864) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9957) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8837);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9441);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9560) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10202) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9932));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10142} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9592} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9970};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10187} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9258} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9266};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8916} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9162} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9925};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9326} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9355} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9662};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8693} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9543} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8762};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9917} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9730} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8938};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10092} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8930} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9116};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9442) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10059} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10136} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9148};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8800, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10140} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10029} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9042} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9625};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9204) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9894) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8966} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8893} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9531};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9559, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9169} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9815} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8670} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9394};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914} = {1'B0, N22225} + {1'B0, N22227} + {1'B0, N22229};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[22], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[21]} = {1'B0, N22040} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9291} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9646};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6231 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6287 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6465 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5959 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6429 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5929 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6242 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[4] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5953 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382} = {1'B0, N21883} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[22]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[22]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8824) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9734) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9954} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9695} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8959};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9376));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8634) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5978 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5985 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6019 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6344 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5960 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6156 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6330 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5972 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6011 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5887 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5912 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6258 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6318 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[1] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6195 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5926 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9505) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9876} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9779} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8783};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8835, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10176} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9080} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9852} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9663};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9271) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9038) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9953) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10129} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8630} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9138};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9597, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9205} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8868} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8695} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9434};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930} = {1'B0, N22241} + {1'B0, N22243} + {1'B0, N22245};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[21], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[20]} = {1'B0, N22048} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8615} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8914};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6501;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6575 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6133 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6030);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6129 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6334 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6091 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[3] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6508 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6008 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104} = {1'B0, N21853} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[21]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[21]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8883) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9573) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9102) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10122} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9589} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9770};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6372 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6297 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5931 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5999 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6174 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6526 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5906 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6059 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6107 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6163 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[0] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6040 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9272)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8994));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8681) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9101} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8756} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9393};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9633, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9887} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8904} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8725};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9799) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9338) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10015) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9945} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8625} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8773};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8673, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9999} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9670} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9472} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10209};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966} = {1'B0, N22314} + {1'B0, N22316} + {1'B0, N22318};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[20], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[19]} = {1'B0, N22056} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8645} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9930};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6087 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6060 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6322 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5973 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6164 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6492 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6273) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6349));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6374 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6450 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6177 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5925 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[2] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6362 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6555 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833} = {1'B0, N21873} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[20]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[20]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8895 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8654));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8735) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8605} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10078} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9006};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8948) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9640) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9172) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9761} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9196} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9387};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10035} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9704} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9507} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8730};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9861) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9403) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10071) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9577} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9939} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10116};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9052} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9480} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10238} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9280};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9402, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9017} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8703} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9244} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9443};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[19], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18]} = {1'B0, N22258} + {1'B0, N22260} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9966};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6542 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6148 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6528 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6010 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6422 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6432 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5992 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6027 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[1] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6204 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6403 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183} = {1'B0, N21863} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[19]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[19]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6484 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6298 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6132 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6378 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6556 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6504 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6402 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6064) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6544 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5911));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6570 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5989) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5962));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[0] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6052 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6554) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N6252 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[22]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10019) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10107) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9924) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9023} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9825} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8876};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10024} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9522} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8589};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9685} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8945} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8890};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9973));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8792) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10072} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10098} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8666};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9007) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9700) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9239) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9377} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8823} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9001};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10214, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9517} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9318} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8583};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9922) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9473) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10134) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9187} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9568} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9755};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9253, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8873} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9288} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10064} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9089};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821} = {1'B0, N22322} + {1'B0, N22324} + {1'B0, N22326};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[18], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]} = {1'B0, N22306} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10182} + {1'B0, N22310};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910} = {1'B0, N22278} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[18]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10171) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10177);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10074) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8827} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8676} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9450};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10144} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8888} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9658};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9037} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9293} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9878};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9605));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8853) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8715} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9712} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9989};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9765) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9982) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8996} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8747} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9178};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9096} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9126} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9865};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9301) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9069) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9536) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10165} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8659} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8816};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9477);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9396) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10229) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9785));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9993} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9810} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10003};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9816));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9984) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10218} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9303} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9786};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9171} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8690} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9105};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9213));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8913) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9812} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10046} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9622};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8838);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9881) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10196) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10232));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9367} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9458} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8736};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8880} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9893} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9650};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10005, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9642} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10043} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9859} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9060};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]} = {1'B0, N22268} + {1'B0, N22270} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9821};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9890) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9202) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8623} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9975} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9423};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10102) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9437) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9672) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9614} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10149} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9798};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9065} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9593} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8643};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10220} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9985} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9259};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9635) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9723) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10044) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10086));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9604) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10045) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10138) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10199) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9436);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10105) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9035} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8707} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9485};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9059} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9863} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9968};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9044);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9514);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9235) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8593) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9626));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9846} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10020} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10041};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10167) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10227) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8696);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10030);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7904);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9073) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8616) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7390));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[2]} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10226} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10067};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9265} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8734} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9791};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9094} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10234} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9339};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8898} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9599} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9665};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8925} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9692} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8987};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10056} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8802} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9076};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8976) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9934} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9428} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9229};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10156} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8809} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8831};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9132) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9826) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9368) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8655} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9807} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9981};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10195} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9227} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9490};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9829, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8910} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9678} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8682};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[15], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[14]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8710} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9421} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9453};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]} = {1'B0, N22286} + {1'B0, N22288} + {1'B0, N22290};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223) | (N22034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8844);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9033) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10081} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9561} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8858};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9268) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9949) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9501) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9606} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9032} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9222};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8952} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10169} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9719};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9838} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8854} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9361};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[14], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9004} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10014} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9030};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307 = !(N22294 & N22296);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10184);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9334} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8721} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10148};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9732) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9414} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9848} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8618};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9198} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8743} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9961};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9619} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10106} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8665};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12028 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9796) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9569) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9168) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8647} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8621} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9840};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8851} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9026} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9754};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8705);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9567) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10010) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9938));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9822));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9099) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9335) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10198} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9214} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8687};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8862} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9629} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9332};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8978} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9494} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9748};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12391 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[12] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9636) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9400) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9860) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10017} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10191} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8679};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9465} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8775} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10204};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10079} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8671} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9100};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9446);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9233) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9273} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9563} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9461};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9471) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9698) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10000} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9653} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9831};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8697} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9369} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9439};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9237} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9530} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9995};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9054);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9298) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8960} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8804} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9068};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9483);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9404) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9918) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9789));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10007} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10089} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10033};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10179} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10115} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9137};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9762) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9534) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8704);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9365) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9405} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9787} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8716};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9263} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9456} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8808};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9110} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9046} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9817};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9601) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8586);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9246) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9823) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9634));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9853} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8882} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9062};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9725} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9570} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8749};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10037);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N7570 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9664);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9433) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9492} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9014} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10051};
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10001} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10151} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9177};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9673);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9998} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9696};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9669) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10222} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10211} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9638};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9331);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9082) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9729) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9474));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9498) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9687} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9871} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9855};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9281);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9565) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9240} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9295};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9147 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8905);
assign {DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2], DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[1]} = {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10207} + {1'B0, DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[19]};
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N10240 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8599);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[1] = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N8931) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9632) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N9310));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[1] & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12155) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12201)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[2]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[2]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[3] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12037 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12433) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12295);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12075) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11879)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[4]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[4]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[5] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12269 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12353) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12213);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11993) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12025)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[6]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[6]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[7] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12340 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12272) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12130);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11916) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12011)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[8]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[8]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[9] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12241 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12191) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12051);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11840) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11847)) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[10]) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[10]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[11] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12134 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11986 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12112) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11974);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203 = ((!N22205) & (!N22199)) | ((!N22201) & (!N22203));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11893 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[13] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169 = !(N22294 | N22296);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425 = (N22194 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12169;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388 = !(((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12307 & N22091) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12203) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12425);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12443) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12388);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445 = !(N22034 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[16] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12445 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12223) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12087);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[17] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[18] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11910);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12368 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12145) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12005);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12305) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12365)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12221);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12254 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11900;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12044 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12183);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12082 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12419) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12283;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12322 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11833);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11965 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12104);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12238 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12382);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11886 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12019);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12160 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12299);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12435 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11943);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12079 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12215);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12358 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11864);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11995 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12137);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12276 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12413);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11921 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12055);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12193 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12335);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11844 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11976);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12116 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12251);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12393 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11897);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12032 | N21818);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12327 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12449 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12311);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838) | N21559;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12091 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11953);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12370 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12225);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12007 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11873);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12287 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12147);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12162 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436 & N20872) | N20876;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11931 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12422);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12204 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12066);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12344 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11853);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11983 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12122);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12178);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12262 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12399);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12042 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11904);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12034 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12004 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12090) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11954;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12144) | N20654;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12199) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12057;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11869 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11977;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023 = N21570 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136 = N21060 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926 = N19751 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12316;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12396;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11850;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12343 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12121) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11980;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12257 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12038) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11903;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12175 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888 = (N21559 & N21570) | N21574;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888 & N21060) | N21064;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12253) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12117;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12367 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11843 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12448) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12310;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050 & N19751) | N19755;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11926) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12417;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[48] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11846) ^ N19431;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[48] & N19158);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18865;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12056;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12218;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12222 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12334;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863 = N21306 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12383;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11911;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280 = N20628 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12070;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12228;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12314) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12174;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12097 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12150) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12012;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11934 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11988) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11856;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12405 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11836) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12325;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12243 & N21306) | N21310;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12081 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12138) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12000;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11923 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11979) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11848;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12086 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12194 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12172) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12031;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410 & N20628) | N20632;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12280) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12141;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12234 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12341 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12200));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[47] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12196 ^ N20265;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[47]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12416;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11944;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11950 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12054;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12105;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12267;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001 = N20621 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12427;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11956;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12035) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11901;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12452 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11876) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12373;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12291 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12348) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12208;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12126 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12184) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12047;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11967 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12023) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11888;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12439 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11865) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12360;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12278 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12336) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12198;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12444 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11920 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11896) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12394;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129 & N20621) | N20625;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12001) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11866;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11829 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12059 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11928));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[46] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11922 ^ N20290;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[46]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12306 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12414;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12103;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363 = N20609 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12426;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12288 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12265) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12125;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11964 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11942) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12436;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12168 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12275 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12250) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12115;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859 & N20609) | N20613;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12363) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12219;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12040 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12418 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12281));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[45] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12277 ^ N20285;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[45]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027 = N20912 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12136;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11834;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12149;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12010 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11987) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11854;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12321 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12298) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12159;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11997 & N20912) | N20916;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12027) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11892;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12083) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11947;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12259 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12142 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12002));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[44] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11999 ^ N20275;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[44]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390 = N20899 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11863;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12182;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12347) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12207;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12045 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12021) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11885;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12357 & N20899) | N20903;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12390) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12246;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12440) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12301;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11852 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11867 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12364));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[43] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12359 ^ N20260;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[43]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111 = N20886 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12216;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11909;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12068) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11933;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12403 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12381) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12239;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12078 & N20886) | N20890;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12111) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11973;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12165) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12024;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12063 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12220 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12084));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[42] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12080 ^ N20280;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[42]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12154;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12016 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11839) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12329;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11889) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12386;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12285 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11948 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12442));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[41] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12438 ^ N20270;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[41]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11881;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12376 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12190) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12050;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12065 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12244) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12106;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11872 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12303 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12166));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[40] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12161 ^ N20295;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[40]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12235;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12100 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11915) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12410;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12372 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11969) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11837;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12089 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12026 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11890));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[39] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11887 ^ N20355;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[39]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11960;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11830 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12271) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12129;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12092 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12326) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12187;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12309 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12387 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12245));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[38] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12242 ^ N20382;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[38]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12318;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12177 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11992) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11859;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12255 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12048) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11912;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11895 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12108 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11971));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[37] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11966 ^ N20370;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[37]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12041;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11906 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12352) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12212;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12407) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12268;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11838 & (!N21559));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[36] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12323 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12114;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[36]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12074) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11937);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12188 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12049));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[35] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12061) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12333;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[35]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12432) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12294);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11913 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12408));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[34] = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11930) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11919;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[34]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12270 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12127));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[33] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12072 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12133;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[33]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11990 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11858));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[32] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12429 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12356;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[32]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12350 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12210));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[31] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12151 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11941;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[31]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12073 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11935));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[30] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11878 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12158;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[30]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12430 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12293));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[29] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12231 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12380;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[29]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12152 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12014));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[28] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11957 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11963;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[28]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13289) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13349)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13325);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13292 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13344) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13285);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11880 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12374));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[27] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12261 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12181;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[27]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12232 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12099));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[26] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11982 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12402;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[26]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13309;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13335 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13293) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13287);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13337 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13318));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13279;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13297 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13345) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13313);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13305 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13330);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13303 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13286));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13329) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13311 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13321);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13277) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13312);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11958 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11827));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[25] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N12345 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N11985;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0] = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[49] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[25]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13278) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13314);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13322) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13340);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13331) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13343)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13275);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13347) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13281);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13290) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13306);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13300) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13284)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13326);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13317 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13294) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13272);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13315) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13333);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20] | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13342) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21])) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13336);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13308) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13270)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13296));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548 = ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13298) & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324)) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13332);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13413) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13324;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13408 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N551;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13410 ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N550;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0] = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N548;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0] ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N549;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[22]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13430 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13478 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13428 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483 = !DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13529 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N683;
assign x[22] = (N22962 & N18245) | ((!N22962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N739);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[11]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[10]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[13]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[12]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[7]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[6]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[9]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[19]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[18]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[21]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13550 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[15]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[14]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[17]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[16]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13449 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13548 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[3]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[2]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[5]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493 = (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[1]) | ((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[0]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13496 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N682;
assign x[21] = (N22964 & N18245) | ((!N22964) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N738);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13486 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13555 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13509 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13573 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13450 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13515 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13465 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13536 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13566 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13514 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13527 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13441 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13577 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13460 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N681;
assign x[20] = (N22966 & N18245) | ((!N22966) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N737);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13456 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13521 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13472 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13542 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13567 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13479 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13435 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13503 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13534 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13477 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13493 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13547) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13561 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13429 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N680;
assign x[19] = (N22965 & N18245) | ((!N22965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N736);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13541 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13559 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13501 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13520 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13448 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13576);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13549 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N679;
assign x[18] = (N22963 & N18245) | ((!N22963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N735);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13508 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13525 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13464 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13485 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13565 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13512);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13516 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N678;
assign x[17] = (N22964 & N18245) | ((!N22964) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N734);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13471 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13492 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13434 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13455 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13533 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13445);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13480 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N677;
assign x[16] = (N22963 & N18245) | ((!N22963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N733);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13440 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13459 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13554 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13572 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13504));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13500 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13451);
assign x[15] = (N22965 & N18245) | ((!N22965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N732);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13507 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13463 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13568);
assign x[14] = (N22965 & N18245) | ((!N22965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N731);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13470 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13433 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13535);
assign x[13] = (N22964 & N18245) | ((!N22964) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N730);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13439 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13553 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13502);
assign x[12] = (N22962 & N18245) | ((!N22962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N729);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13491 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13519 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13466);
assign x[11] = (N22962 & N18245) | ((!N22962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N728);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13546 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13484 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13436);
assign x[10] = (N22964 & N18245) | ((!N22964) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N727);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13444 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13454 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13556);
assign x[9] = (N22966 & N18245) | ((!N22966) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N726);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13498 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13571 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13522);
assign x[8] = (N22965 & N18245) | ((!N22965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N725);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874 = !((DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13540 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N18874);
assign x[7] = (N22962 & N18245) | ((!N22962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N724);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13543);
assign x[6] = (N22963 & N18245) | ((!N22963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N723);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13473);
assign x[5] = (N22963 & N18245) | ((!N22963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N722);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13560);
assign x[4] = (N22963 & N18245) | ((!N22963) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N721);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13494);
assign x[3] = (N22965 & N18245) | ((!N22965) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N720);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13578);
assign x[2] = (N22966 & N18245) | ((!N22966) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N719);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13513);
assign x[1] = (N22964 & N18245) | ((!N22964) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N718);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717 = !(((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13483) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13447);
assign x[0] = (N22962 & N18245) | ((!N22962) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N717);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585 = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__68 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N494;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N585 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82));
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[30] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13897 & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N595;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13469));
assign x[27] = (N18402 & N18406) | ((!N18402) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N713);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13489));
assign x[26] = (N18402 & N18406) | ((!N18402) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N712);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13487));
assign x[25] = (N18402 & N18406) | ((!N18402) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N711);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13532));
assign x[24] = (N18402 & N18406) | ((!N18402) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N710);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13757 & (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13539));
assign x[23] = (N18402 & N18406) | ((!N18402) & DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N709);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[6] | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__82);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708 = !(DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N5563 | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[4]);
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493 = (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N708) ^ DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N707;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[31] = !((((!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N13872) | (!DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_N493)) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[8]) | DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[7]);
reg x_reg_28__I3792_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I3792_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29];
	end
assign x[28] = x_reg_28__I3792_QOUT;
reg x_reg_30__I3794_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I3794_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[30];
	end
assign x[30] = x_reg_30__I3794_QOUT;
reg x_reg_31__I3795_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I3795_QOUT <= DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[31];
	end
assign x[31] = x_reg_31__I3795_QOUT;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[28] = DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[29];
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__42[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__61[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__195[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[1] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[2] = 1'B0;
assign DFT_compute_cynw_cm_float_cos_E8_M23_2_inst_inst_cellmath__215[4] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urP3TQjXoxlO : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



