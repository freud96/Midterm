/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:55 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195;
wire [20:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197;
wire [32:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122,
	DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129;
wire N19976,N19980,N19983,N19994,N19998,N20199,N20253 
	,N20260,N20350,N20360,N20370,N20392,N20414,N20424,N20434 
	,N20444,N20454,N20471,N20481,N20491,N20501,N20537,N20547 
	,N20557,N20567,N20577,N20587,N20597,N20607,N20617,N20988 
	,N21042,N21116,N21208,N21231,N21450,N21461,N21468,N21766 
	,N21801,N22304,N22319,N22330,N22332,N22342,N22344,N22349 
	,N22351,N22356,N22358,N22361,N22366,N22368,N22373,N22378 
	,N22385,N22387,N22392,N22395,N22397,N22402,N22404,N22409 
	,N22411,N22416,N22421,N22423,N22430,N22432,N22437,N22439 
	,N22442,N22444,N22451,N22453,N22482,N22484,N22489,N22504 
	,N22508,N22510,N22512,N22516,N22518,N22520,N22524,N22526 
	,N22528,N22531,N22534,N22536,N22558,N22562,N22564,N22566 
	,N22569,N22571,N22581,N22583,N22593,N22598,N22600,N22644 
	,N22646,N22648,N23029,N23056,N23313,N23314,N23315,N23316 
	,N23317,N23318,N23319,N23320,N23321,N23322,N23323,N23324 
	,N23325,N23326,N23327,N23328,N23329,N23330,N23331,N23332 
	,N23333,N23334,N23335,N23336;
reg x_reg_31__retimed_I13794_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13794_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990;
	end
assign N23056 = x_reg_31__retimed_I13794_QOUT;
reg x_reg_31__retimed_I13781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13781_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441;
	end
assign N23029 = x_reg_31__retimed_I13781_QOUT;
reg x_reg_31__retimed_I13653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13653_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700;
	end
assign N22648 = x_reg_31__retimed_I13653_QOUT;
reg x_reg_31__retimed_I13652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13652_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649;
	end
assign N22646 = x_reg_31__retimed_I13652_QOUT;
reg x_reg_31__retimed_I13651_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13651_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896;
	end
assign N22644 = x_reg_31__retimed_I13651_QOUT;
reg x_reg_31__retimed_I13631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13631_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089;
	end
assign N22600 = x_reg_31__retimed_I13631_QOUT;
reg x_reg_31__retimed_I13630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13630_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959;
	end
assign N22598 = x_reg_31__retimed_I13630_QOUT;
reg x_reg_31__retimed_I13628_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13628_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822;
	end
assign N22593 = x_reg_31__retimed_I13628_QOUT;
reg x_reg_31__retimed_I13625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13625_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015;
	end
assign N22583 = x_reg_31__retimed_I13625_QOUT;
reg x_reg_31__retimed_I13624_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13624_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888;
	end
assign N22581 = x_reg_31__retimed_I13624_QOUT;
reg x_reg_31__retimed_I13620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13620_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761;
	end
assign N22571 = x_reg_31__retimed_I13620_QOUT;
reg x_reg_31__retimed_I13619_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13619_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644;
	end
assign N22569 = x_reg_31__retimed_I13619_QOUT;
reg x_reg_31__retimed_I13618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13618_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783;
	end
assign N22566 = x_reg_31__retimed_I13618_QOUT;
reg x_reg_31__retimed_I13617_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13617_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028;
	end
assign N22564 = x_reg_31__retimed_I13617_QOUT;
reg x_reg_31__retimed_I13616_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13616_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911;
	end
assign N22562 = x_reg_31__retimed_I13616_QOUT;
reg x_reg_31__retimed_I13615_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13615_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830;
	end
assign N22558 = x_reg_31__retimed_I13615_QOUT;
reg x_reg_31__retimed_I13608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13608_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655;
	end
assign N22536 = x_reg_31__retimed_I13608_QOUT;
reg x_reg_31__retimed_I13607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13607_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006;
	end
assign N22534 = x_reg_31__retimed_I13607_QOUT;
reg x_reg_31__retimed_I13606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13606_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634;
	end
assign N22531 = x_reg_31__retimed_I13606_QOUT;
reg x_reg_31__retimed_I13605_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13605_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712;
	end
assign N22528 = x_reg_31__retimed_I13605_QOUT;
reg x_reg_31__retimed_I13604_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13604_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861;
	end
assign N22526 = x_reg_31__retimed_I13604_QOUT;
reg x_reg_31__retimed_I13603_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13603_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841;
	end
assign N22524 = x_reg_31__retimed_I13603_QOUT;
reg x_reg_31__retimed_I13602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13602_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537;
	end
assign N22520 = x_reg_31__retimed_I13602_QOUT;
reg x_reg_31__retimed_I13601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13601_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666;
	end
assign N22518 = x_reg_31__retimed_I13601_QOUT;
reg x_reg_31__retimed_I13600_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13600_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902;
	end
assign N22516 = x_reg_31__retimed_I13600_QOUT;
reg x_reg_31__retimed_I13599_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13599_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039;
	end
assign N22512 = x_reg_31__retimed_I13599_QOUT;
reg x_reg_31__retimed_I13598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13598_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610;
	end
assign N22510 = x_reg_31__retimed_I13598_QOUT;
reg x_reg_31__retimed_I13597_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13597_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590;
	end
assign N22508 = x_reg_31__retimed_I13597_QOUT;
reg x_reg_31__retimed_I13596_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13596_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951;
	end
assign N22504 = x_reg_31__retimed_I13596_QOUT;
reg x_reg_31__retimed_I13591_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13591_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787;
	end
assign N22489 = x_reg_31__retimed_I13591_QOUT;
reg x_reg_31__retimed_I13589_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13589_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980;
	end
assign N22484 = x_reg_31__retimed_I13589_QOUT;
reg x_reg_31__retimed_I13588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13588_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859;
	end
assign N22482 = x_reg_31__retimed_I13588_QOUT;
reg x_reg_31__retimed_I13586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13586_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014;
	end
assign N22453 = x_reg_31__retimed_I13586_QOUT;
reg x_reg_31__retimed_I13585_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13585_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564;
	end
assign N22451 = x_reg_31__retimed_I13585_QOUT;
reg x_reg_31__retimed_I13582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13582_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652;
	end
assign N22444 = x_reg_31__retimed_I13582_QOUT;
reg x_reg_31__retimed_I13581_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13581_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525;
	end
assign N22442 = x_reg_31__retimed_I13581_QOUT;
reg x_reg_31__retimed_I13580_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13580_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619;
	end
assign N22439 = x_reg_31__retimed_I13580_QOUT;
reg x_reg_31__retimed_I13579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13579_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739;
	end
assign N22437 = x_reg_31__retimed_I13579_QOUT;
reg x_reg_31__retimed_I13577_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13577_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877;
	end
assign N22432 = x_reg_31__retimed_I13577_QOUT;
reg x_reg_31__retimed_I13576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13576_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000;
	end
assign N22430 = x_reg_31__retimed_I13576_QOUT;
reg x_reg_31__retimed_I13573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13573_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024;
	end
assign N22423 = x_reg_31__retimed_I13573_QOUT;
reg x_reg_31__retimed_I13572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13572_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899;
	end
assign N22421 = x_reg_31__retimed_I13572_QOUT;
reg x_reg_31__retimed_I13570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13570_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571;
	end
assign N22416 = x_reg_31__retimed_I13570_QOUT;
reg x_reg_31__retimed_I13568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13568_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958;
	end
assign N22411 = x_reg_31__retimed_I13568_QOUT;
reg x_reg_31__retimed_I13567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13567_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840;
	end
assign N22409 = x_reg_31__retimed_I13567_QOUT;
reg x_reg_31__retimed_I13565_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13565_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589;
	end
assign N22404 = x_reg_31__retimed_I13565_QOUT;
reg x_reg_31__retimed_I13564_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13564_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038;
	end
assign N22402 = x_reg_31__retimed_I13564_QOUT;
reg x_reg_31__retimed_I13562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13562_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782;
	end
assign N22397 = x_reg_31__retimed_I13562_QOUT;
reg x_reg_31__retimed_I13561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13561_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665;
	end
assign N22395 = x_reg_31__retimed_I13561_QOUT;
reg x_reg_31__retimed_I13560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13560_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669;
	end
assign N22392 = x_reg_31__retimed_I13560_QOUT;
reg x_reg_31__retimed_I13558_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13558_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703;
	end
assign N22387 = x_reg_31__retimed_I13558_QOUT;
reg x_reg_31__retimed_I13557_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13557_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826;
	end
assign N22385 = x_reg_31__retimed_I13557_QOUT;
reg x_reg_31__retimed_I13554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13554_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964;
	end
assign N22378 = x_reg_31__retimed_I13554_QOUT;
reg x_reg_31__retimed_I13552_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13552_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811;
	end
assign N22373 = x_reg_31__retimed_I13552_QOUT;
reg x_reg_31__retimed_I13550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13550_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760;
	end
assign N22368 = x_reg_31__retimed_I13550_QOUT;
reg x_reg_31__retimed_I13549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13549_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643;
	end
assign N22366 = x_reg_31__retimed_I13549_QOUT;
reg x_reg_31__retimed_I13547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13547_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528;
	end
assign N22361 = x_reg_31__retimed_I13547_QOUT;
reg x_reg_31__retimed_I13546_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13546_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079;
	end
assign N22358 = x_reg_31__retimed_I13546_QOUT;
reg x_reg_31__retimed_I13545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13545_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630;
	end
assign N22356 = x_reg_31__retimed_I13545_QOUT;
reg x_reg_31__retimed_I13543_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13543_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804;
	end
assign N22351 = x_reg_31__retimed_I13543_QOUT;
reg x_reg_31__retimed_I13542_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13542_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800;
	end
assign N22349 = x_reg_31__retimed_I13542_QOUT;
reg x_reg_31__retimed_I13540_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13540_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061;
	end
assign N22344 = x_reg_31__retimed_I13540_QOUT;
reg x_reg_31__retimed_I13539_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13539_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609;
	end
assign N22342 = x_reg_31__retimed_I13539_QOUT;
reg x_reg_31__retimed_I13535_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13535_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432;
	end
assign N22332 = x_reg_31__retimed_I13535_QOUT;
reg x_reg_31__retimed_I13534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13534_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446;
	end
assign N22330 = x_reg_31__retimed_I13534_QOUT;
reg x_reg_31__retimed_I13531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13531_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881;
	end
assign N22319 = x_reg_31__retimed_I13531_QOUT;
reg x_reg_31__retimed_I13526_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13526_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614;
	end
assign N22304 = x_reg_31__retimed_I13526_QOUT;
reg x_reg_31__retimed_I13362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13362_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543;
	end
assign N21801 = x_reg_31__retimed_I13362_QOUT;
reg x_reg_31__retimed_I13349_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13349_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22];
	end
assign N21766 = x_reg_31__retimed_I13349_QOUT;
reg x_reg_31__retimed_I13270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13270_QOUT <= a_exp[5];
	end
assign N21468 = x_reg_31__retimed_I13270_QOUT;
reg x_reg_31__retimed_I13267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13267_QOUT <= a_exp[6];
	end
assign N21461 = x_reg_31__retimed_I13267_QOUT;
reg x_reg_31__retimed_I13262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13262_QOUT <= a_exp[0];
	end
assign N21450 = x_reg_31__retimed_I13262_QOUT;
reg x_reg_31__retimed_I13187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13187_QOUT <= a_exp[2];
	end
assign N21231 = x_reg_31__retimed_I13187_QOUT;
reg x_reg_31__retimed_I13177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13177_QOUT <= a_exp[1];
	end
assign N21208 = x_reg_31__retimed_I13177_QOUT;
reg x_reg_31__retimed_I13151_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13151_QOUT <= a_exp[3];
	end
assign N21116 = x_reg_31__retimed_I13151_QOUT;
reg x_reg_31__retimed_I13120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13120_QOUT <= a_exp[4];
	end
assign N21042 = x_reg_31__retimed_I13120_QOUT;
reg x_reg_31__retimed_I13108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I13108_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647;
	end
assign N20988 = x_reg_31__retimed_I13108_QOUT;
reg x_reg_31__retimed_I12961_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12961_QOUT <= a_man[0];
	end
assign N20617 = x_reg_31__retimed_I12961_QOUT;
reg x_reg_31__retimed_I12957_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12957_QOUT <= a_man[1];
	end
assign N20607 = x_reg_31__retimed_I12957_QOUT;
reg x_reg_31__retimed_I12953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12953_QOUT <= a_man[2];
	end
assign N20597 = x_reg_31__retimed_I12953_QOUT;
reg x_reg_31__retimed_I12949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12949_QOUT <= a_man[8];
	end
assign N20587 = x_reg_31__retimed_I12949_QOUT;
reg x_reg_31__retimed_I12945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12945_QOUT <= a_man[7];
	end
assign N20577 = x_reg_31__retimed_I12945_QOUT;
reg x_reg_31__retimed_I12941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12941_QOUT <= a_man[4];
	end
assign N20567 = x_reg_31__retimed_I12941_QOUT;
reg x_reg_31__retimed_I12937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12937_QOUT <= a_man[15];
	end
assign N20557 = x_reg_31__retimed_I12937_QOUT;
reg x_reg_31__retimed_I12933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12933_QOUT <= a_man[21];
	end
assign N20547 = x_reg_31__retimed_I12933_QOUT;
reg x_reg_31__retimed_I12929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12929_QOUT <= a_man[17];
	end
assign N20537 = x_reg_31__retimed_I12929_QOUT;
reg x_reg_31__retimed_I12914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12914_QOUT <= a_man[3];
	end
assign N20501 = x_reg_31__retimed_I12914_QOUT;
reg x_reg_31__retimed_I12910_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12910_QOUT <= a_man[5];
	end
assign N20491 = x_reg_31__retimed_I12910_QOUT;
reg x_reg_31__retimed_I12906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12906_QOUT <= a_man[11];
	end
assign N20481 = x_reg_31__retimed_I12906_QOUT;
reg x_reg_31__retimed_I12902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12902_QOUT <= a_man[10];
	end
assign N20471 = x_reg_31__retimed_I12902_QOUT;
reg x_reg_31__retimed_I12895_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12895_QOUT <= a_man[19];
	end
assign N20454 = x_reg_31__retimed_I12895_QOUT;
reg x_reg_31__retimed_I12891_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12891_QOUT <= a_man[16];
	end
assign N20444 = x_reg_31__retimed_I12891_QOUT;
reg x_reg_31__retimed_I12887_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12887_QOUT <= a_man[12];
	end
assign N20434 = x_reg_31__retimed_I12887_QOUT;
reg x_reg_31__retimed_I12883_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12883_QOUT <= a_man[9];
	end
assign N20424 = x_reg_31__retimed_I12883_QOUT;
reg x_reg_31__retimed_I12879_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12879_QOUT <= a_man[14];
	end
assign N20414 = x_reg_31__retimed_I12879_QOUT;
reg x_reg_31__retimed_I12870_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12870_QOUT <= a_man[20];
	end
assign N20392 = x_reg_31__retimed_I12870_QOUT;
reg x_reg_31__retimed_I12861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12861_QOUT <= a_man[6];
	end
assign N20370 = x_reg_31__retimed_I12861_QOUT;
reg x_reg_31__retimed_I12857_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12857_QOUT <= a_man[13];
	end
assign N20360 = x_reg_31__retimed_I12857_QOUT;
reg x_reg_31__retimed_I12853_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12853_QOUT <= a_man[18];
	end
assign N20350 = x_reg_31__retimed_I12853_QOUT;
reg x_reg_22__retimed_I12816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12816_QOUT <= a_man[22];
	end
assign N20260 = x_reg_22__retimed_I12816_QOUT;
reg x_reg_31__retimed_I12813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12813_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612;
	end
assign N20253 = x_reg_31__retimed_I12813_QOUT;
reg x_reg_26__retimed_I12789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__retimed_I12789_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580;
	end
assign N20199 = x_reg_26__retimed_I12789_QOUT;
reg x_reg_22__retimed_I12700_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12700_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759;
	end
assign N19998 = x_reg_22__retimed_I12700_QOUT;
assign N23313 = !N19998;
assign N23319 = !N23313;
assign N23318 = !N23313;
assign N23317 = !N23313;
assign N23316 = !N23313;
assign N23315 = !N23313;
assign N23314 = !N23313;
reg x_reg_22__retimed_I12698_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I12698_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646;
	end
assign N19994 = x_reg_22__retimed_I12698_QOUT;
assign N23320 = !N19994;
assign N23326 = !N23320;
assign N23325 = !N23320;
assign N23324 = !N23320;
assign N23323 = !N23320;
assign N23322 = !N23320;
assign N23321 = !N23320;
reg x_reg_20__retimed_I12693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I12693_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82;
	end
assign N19983 = x_reg_20__retimed_I12693_QOUT;
assign N23327 = !N19983;
assign N23328 = !N23327;
reg x_reg_31__retimed_I12692_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12692_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639;
	end
assign N19980 = x_reg_31__retimed_I12692_QOUT;
assign N23329 = !N19980;
assign N23336 = !N23329;
assign N23335 = !N23329;
assign N23334 = !N23329;
assign N23333 = !N23329;
assign N23332 = !N23329;
assign N23331 = !N23329;
assign N23330 = !N23329;
reg x_reg_31__retimed_I12690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I12690_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829;
	end
assign N19976 = x_reg_31__retimed_I12690_QOUT;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746 = !(a_exp[6] & a_exp[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749 = !(a_exp[4] & a_exp[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737 = !(a_exp[2] & a_exp[1]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738 = !((a_exp[7] & a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15744);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15746 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22738);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15854;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839 = !(a_sign & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829 = !a_sign;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__19);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798 = !(a_man[4] | a_man[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15798 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15767) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15777) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15788;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956 = !a_man[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790 = !(a_man[0] | a_man[1]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15790);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053 = !(a_man[22] | a_man[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763 = !(a_man[20] | a_man[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804 = !(a_man[12] | a_man[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773 = !(a_man[18] | a_man[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784 = !(a_man[16] | a_man[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794 = !(a_man[14] | a_man[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15804 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15773) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15784) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15794;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15763) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15796);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15771 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22746);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15780 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15769);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15832 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15839) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__24);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863 = ((a_exp[7] | a_exp[6]) | a_exp[0]) | a_exp[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867 = ((a_exp[4] | a_exp[2]) | a_exp[3]) | a_exp[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15863 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15867);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__17 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__68) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898 = !(a_exp[5] & a_exp[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15898);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639 = !(a_exp[7] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15891);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100 = !a_exp[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103 = !a_exp[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107 = !a_exp[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070 = !(a_exp[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 = (!a_exp[5]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44070;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7107 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7108;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] = a_exp[4] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7102;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236 = !(a_man[22] & a_man[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190 = !a_man[21];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177} = {1'B0, a_man[20]} + {1'B0, a_man[22]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802} = {1'B0, a_man[19]} + {1'B0, a_man[21]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816 = !a_man[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454 = a_man[12] | a_man[14];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816} + {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5454};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912 = (!a_man[14]) ^ a_man[16];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211 = a_man[13] | a_man[15];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587} = {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6211};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5912} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5406} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5587};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798 = (!a_man[15]) ^ a_man[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103 = a_man[14] | a_man[16];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703 = !a_man[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966} = {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6103} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5798} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5773} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5966};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437 = !a_man[19];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748} = {1'B0, a_man[11]} + {1'B0, a_man[13]} + {1'B0, a_man[16]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699} = {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5944};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028 = (!a_man[13]) ^ a_man[15];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6028} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5887} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6083};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541 = !a_man[17];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926 = !a_man[18];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862} = {1'B0, a_man[10]} + {1'B0, a_man[12]} + {1'B0, a_man[15]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5558} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6059};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132 = (!a_man[12]) ^ a_man[14];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6132} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5507} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5699};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975} = {1'B0, a_man[9]} + {1'B0, a_man[11]} + {1'B0, a_man[14]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6163} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6243} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5862};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5748} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6185} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6004};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854} = {1'B0, a_man[17]} + {1'B0, a_man[19]} + {1'B0, a_man[22]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427} = {1'B0, a_man[18]} + {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6051};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040 = !a_man[16];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476} = {1'B0, a_man[18]} + {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5668} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5854};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992 = a_man[15] | a_man[17];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5992} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5476} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6155};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951 = a_man[22] | a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659 = !a_man[15];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090} = {1'B0, a_man[10]} + {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754 = (!a_man[22]) ^ a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252} = {1'B0, a_man[21]} + {1'B0, a_man[7]} + {1'B0, a_man[9]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5571} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5754} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5414} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5975} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5783};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5676} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5810} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5621};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147 = !a_man[14];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491} = {1'B0, a_man[20]} + {1'B0, a_man[6]} + {1'B0, a_man[8]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761 = !a_man[13];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761} + {1'B0, a_man[11]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6064} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5683} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6252};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5514} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6090} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5895};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5485} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5433} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6115};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399 = !a_man[12];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6173};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605} = {1'B0, a_man[19]} + {1'B0, a_man[5]} + {1'B0, a_man[7]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5872} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5491};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6193} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5627} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6011};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5727} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5921};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878 = !a_man[11];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5421} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715} = {1'B0, a_man[18]} + {1'B0, a_man[4]} + {1'B0, a_man[6]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5985} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5905} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5605};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5736} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5441} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6123};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6221} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5708} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5535};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496 = !a_man[10];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496} + {1'B0, a_man[8]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5522} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852} = {1'B0, a_man[17]} + {1'B0, a_man[3]} + {1'B0, a_man[5]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6021} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6097} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5715};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5847} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5544} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6227};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5818} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5842} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6036};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862} = {1'B0, a_man[16]} + {1'B0, a_man[2]} + {1'B0, a_man[4]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43875};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993 = !a_man[9];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43881} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43837} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43852};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5957} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5661} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5468};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5929} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5460} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5654};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478 = a_man[22] | a_man[15];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054} = {1'B0, a_man[1]} + {1'B0, a_man[3]} + {1'B0, a_man[6]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5478} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6237};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612 = !a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43845} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43862} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43890};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43884} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43841} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43870};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6043} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5953} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6143};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889} = {1'B0, a_man[21]} + {1'B0, a_man[14]} + {1'B0, a_man[0]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105 = !a_man[7];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408} = {1'B0, a_man[2]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6085} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5969} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5590};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156 = (!a_man[22]) ^ a_man[15];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6054} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6156} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43831};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43849} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43894} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43878};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43853} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43846} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43867};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434 = a_man[20] | a_man[13];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760 = !a_man[6];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488} = {1'B0, a_man[1]} + {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5434} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5700} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6188};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5775} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5408} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5889};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43834} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43859} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43887};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43891} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43856} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43838};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473 = (!a_man[20]) ^ a_man[13];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43517} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43473} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43488};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656 = a_man[19] | a_man[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212 = !a_man[5];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481} = {1'B0, a_man[0]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5656} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43526} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43498};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5530} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5914} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6108};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5499} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5685} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5874};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990 = a_man[17] | a_man[10];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5990} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5397};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574} = {1'B0, a_man[18]} + {1'B0, a_man[11]} + {1'B0, a_man[2]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833 = !a_man[4];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5758} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6145};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551 = !a_man[3];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5876} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5574} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5955};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43530} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43485} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43514};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467 = (!a_man[19]) ^ a_man[12];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43467} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43511} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43481};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43506} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43477} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43520};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43489} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43482} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43503};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5614} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6174} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5493};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560 = !a_man[1];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580 = !a_man[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840 = a_man[5] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5840} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5702} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5534} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5890};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919} = {1'B0, a_man[7]} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5726} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5431} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5919} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6086} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5409};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808} = {1'B0, a_man[8]} + {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5620} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6113} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5808};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6183} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5591} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5779};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651 = (!a_man[5]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007} = {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6189} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5651} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5510};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624} = {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878} + {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5436} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5624};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5813} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6007} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5538} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5731} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5924} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6120} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6153;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5577} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6235);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6026 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5467) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6148);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6128);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5448 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5636);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5660 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6226) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6042);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6176) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5398)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6068);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5823 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6019);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5730 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5734) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5542);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5464} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5658} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5845} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6203 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5714 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5904);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5928 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5626) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5439);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5857) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5778)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5671);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6039} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6225};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6010;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6096 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5420);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5603 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5791);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6192;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44036) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5512 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5817);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5606) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5503);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5984 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6172);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5681);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5707 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5413) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6089);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5871 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6063);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6249 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5569);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5594 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6162) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5973);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6050) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5965)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5852));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6081) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5976)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5786);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5753 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5950);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5540 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6121) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5927);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6140 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5459);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5650 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5839);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5438 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6008) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5814);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5936) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6020)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5825);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815 = (!a_man[9]) ^ a_man[2];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5815} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5399};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6001} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5505} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5695};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5970} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6079} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6159};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009 = a_man[9] | a_man[2];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705} = {1'B0, a_man[10]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5705} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6009} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5761};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5585} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5886} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5404};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5481} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5961} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5672};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088} = {1'B0, a_man[11]} + {1'B0, a_man[4]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5891} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6147} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6088};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22553} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5473} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5770} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6152};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5851} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5858} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6056};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592} = {1'B0, a_man[12]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5551};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5659} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5411} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5592};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5664} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6231} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6047};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5740} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6239} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5555};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5410);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5682 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6033 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6218);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5533 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5724);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5893 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6191) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5917 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6111);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5430 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5619);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6087 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5780) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5492) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5570)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6251);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674 = a_man[14] | a_man[7];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5674};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5993};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484 = (!a_man[14]) ^ a_man[7];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972} = {1'B0, a_man[13]} + {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5833};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6212} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5580};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6160} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5484} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6241};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6199} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5900} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5711};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025 = (!a_man[16]) ^ a_man[9];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5703} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5878};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5956} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6105};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5425} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6025} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5909};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941 = a_man[15] | a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5496} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5760} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5560};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5941} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5829};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746 = (!a_man[15]) ^ a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5556} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5746} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5642};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5788} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6093} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5600};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6169} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6023} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6207};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795 = (!a_man[17]) ^ a_man[10];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6066} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5795} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5687};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209 = a_man[16] | a_man[9];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6209} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5610} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6100};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5980} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5488};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6061} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5523} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5718};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43470} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43495} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43523};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5946} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5907} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6098};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43492} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43527} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43474};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5934} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5612};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5549} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6126} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5932};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6040} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5781} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5972};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5445} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6014} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5820};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5517} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5451};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5417} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5640} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5826};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5632} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5744} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5939};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6161 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5806 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6182 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5504);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5971 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5673) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5483);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5693 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5885);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5403 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6078);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6002)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5807);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5583 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5768);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5960 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6151);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5471 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5850 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6046);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5548)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6232);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6230 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5546);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5739 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5931);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6125 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5444);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5819 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5631);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5979)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5789);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6012 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6198);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5516 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5710);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5898 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6091);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5416 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5529)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6214);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5787 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6168 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5486);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5677 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5866);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6245 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6060);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5958)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5764);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5562 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5945 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5455 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5645);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5835 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5513)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6213 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5528);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5721 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5913);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5427 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6107);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5802 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5613);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5943)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5747);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5720) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5526;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5967) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5776);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5794)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5607);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6222) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6035);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5994 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6177);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6190 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5426 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5821)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5633));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6236 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6053));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6038 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5978;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5487 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5844;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6124) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5442));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248 = !(a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1] = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5968 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5774));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6101)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5910);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6210 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6045;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5547 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5576;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6200);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6220);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5604;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6034 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5769) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5584);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6013 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5751) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5564);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5996 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5735) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5543);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5422)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6099);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5841) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5849) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6044));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5589 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5407));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6058;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5863;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5796);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5991 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5694;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6077 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6070;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6150) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5469));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5856 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5684) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5545) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5738));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5477 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6158));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5987) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5588;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[1]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7100) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43412;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7181 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6187 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6006));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5831 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5453)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5521;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5903 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5586;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6181) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5501));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5811 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5623));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5628 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6052;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5552 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5440;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5618) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5805));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6084 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6219;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5725 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5688;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5582) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5701 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5508));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5974;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6165));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5870;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6250 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5962;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5884) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6076));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7213));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7197));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7160);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N752;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N634) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N635));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N636) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N637));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N630) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N631));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N632) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N633));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5435 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6117));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5480) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5916) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6110));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N627));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N628) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N629));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7341 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44063) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7361);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N751;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7248);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7136) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7281));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7168) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7311));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5922 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5729));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5777) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6082;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N626));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7203) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7306);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N750;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7157) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7128));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7330 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N755;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7350 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7357) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7325));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7162));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7273);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N754;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7192);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7335) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7225));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7367) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22759 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7307) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7217);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N753;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7746 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7832);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8162;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[21] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8060);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[18] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8108 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8500 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[22] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8274 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[19] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8130;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8707;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7929 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8745);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8739);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7904);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[29] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7956 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8438) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8288) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7809);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[29];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8290);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8489 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8463;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7941);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8417 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8173);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843 = 1'B0 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8384 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8723);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7689);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8425);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8238) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8484)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8098);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[27] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7867) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8444) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[27]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14655 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5655 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5463));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5812) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5938;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5828) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5906)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5717);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5461) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6142);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5948) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6139));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6144 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5954));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6119) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5536 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6244 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5675)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6116;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6184 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5622;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6216) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5532));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6037 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5843));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6073 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5756;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5880 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6141;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5648) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5698) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5838));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7135));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7304) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7269));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7339);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N746;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N624) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N625));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7147) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5759 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5573));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5784);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5892)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5827;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6205 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5920;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5639);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6157;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5450) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5524)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6206);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5479 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5952) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5757);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N621));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N622) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N623));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7194) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7212));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7184));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7283);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N745;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7289) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7176));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7190));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7324);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7152));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7140);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N747;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12783 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11832 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7807;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8390 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8634);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7881 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8685);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8459 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7827;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7997 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8389;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8663;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8757);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7741);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7954 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8191;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11294) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7346) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5396 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6067));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5646 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5482;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5859 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5457;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5680) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5869));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N620));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7124) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7337) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7156));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7327));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7229);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N744;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5875 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5686));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6146) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5983) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6171));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N619));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7322) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7222));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7227) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7355));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7215));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7173);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N743;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22721;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12814 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11862 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8244 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8492);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8536 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8341);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8493 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7959 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7969 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7712;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8609);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8752)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8225) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8710);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N780;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11192) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5494 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6175));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N618));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7166 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44056) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7171) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7299));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7359));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7371);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22642;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7334) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7301));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5989 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5797));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44043 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5732) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5539;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5925 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5652;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5394;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288 = !a_exp[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7210) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7354));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7365));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7270) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7239));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7245));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7316);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N741;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12844 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11813} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12730} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11562};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7278) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7125);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7263));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N748;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7249) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7252);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N749;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12753 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42] = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11796 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8170;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7923) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7699;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8061)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8632;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8257);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7721 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8517);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7834 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8690;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11327) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12847) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11230) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12199} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11389};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12345} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11623} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11559};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11897 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11162) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5609 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5424));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6092 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6069;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5899 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5578;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N616));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7310));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7315) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7189));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7146) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7138));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7261);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N740;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43262);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245 = !(a_exp[0] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43255);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6102 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5908));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5611;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43261 | (!a_exp[0]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43245) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43242 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6186;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43289 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43236) | a_exp[0]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43285 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43288) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43266);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43268) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43251);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43233 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43271);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7255));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7259) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7134));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7347) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7280));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7206);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N739;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12875 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11259) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12237} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11428};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8414;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8116);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8211));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8305;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8776;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8759);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8497;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8017;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7759;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8313) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8563);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8046 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8419);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8618 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7791 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8525) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7747);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N776;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11390) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11968} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11312} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11246};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8441;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8449);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7964 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8549 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8297);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8256;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7928 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8783;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11461) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11356) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11326) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11226) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11852} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12763} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11625};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12381} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11575} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11214};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8457);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8472);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8637;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7669 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7733);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8571 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7936);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8674));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8032);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8605 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8705);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7986 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7688);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8182 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8424;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11524) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11424) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11189) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43280) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43267));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5719 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5525));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5911) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5554;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7298) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7200));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7204) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7333));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7290) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7224));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7151);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N738;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6208 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6024));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5737 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5579)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44049) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6133) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5643 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6253;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5873;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5447) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5635));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N613));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N614) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N615));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7243) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7144));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7149) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7276));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7169));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7352);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22635;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11186 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11291) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12273} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11467};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12012} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11195} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12840};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12661} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12715} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11683};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12087} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12742} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12805};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[38], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[37]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11398} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12330} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12174};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8736;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8475;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8671);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8366;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8653) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8455) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8120 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8138);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[19] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8511) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7730) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[13];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9945} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9909} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10070};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9992} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10349} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10308};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9960} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9930} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10159};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10489} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10086} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10278};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10416} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10234} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10025};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10384} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10334} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10432};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9937} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10066} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9914};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10208} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10147} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10484};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10046} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10103} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10318};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10413} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10528} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10286};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10263} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10509} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10478};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10012} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10014} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10281};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9908} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10125} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10180};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10140} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10133} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10356};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10149} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10362} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10505};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9995} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10198} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10059};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10170} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10512} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10442};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10338} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9932} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9991};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10498} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10224} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9929};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10328} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10038} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10307};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10150} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10418} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10094};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10214} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10511} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10526};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10342} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9946} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9922};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10078} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10276} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10091};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9942} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10423} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10011};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10226} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3658} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10237};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10182} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10456} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10431};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10191} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10218} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10500};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10245} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9980} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9959};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5830 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5641));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5665 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5785;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5472 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6164;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5935));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N612));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7187) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7121) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7344));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7349) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7220));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7178) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7368));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7293);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N736;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10294} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9970};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9982} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9955} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10419};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5452 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6131));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5942;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6049) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N611));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7132) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7319) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7287));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7292) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7165));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7123) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43414);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43404;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10319} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10306} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9975};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5940 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5745));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6242) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6238;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N610));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7331) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7233));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7364));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7321) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7182);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N734;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22602;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10305} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10521} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10062};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10353} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10386} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10310};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10154} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10024} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10090};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10421} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10439} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10329};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10040} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10284} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9935};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10339} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9971} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9993};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10050} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10075} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10321};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10085} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10104} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10371};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10348} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10029} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10002};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10471} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10136} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10113};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10518} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10049} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10324};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5557 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6057;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5918);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6075 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5860);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6112) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5800)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5986);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N6228) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5848;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5669) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N5475));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163 = !((a_exp[0] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N608) | ((!a_exp[0]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N609));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7275) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7163));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7209) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7271) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7175));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7179) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[4]) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7309));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7267) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7202));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7127);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7631) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N733;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10409} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10168};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10087} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10004} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10271};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10538} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10172} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10247};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10206} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9961} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10228};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10238} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10260} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10527};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10037) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10508;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10054} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10396};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[15]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10126} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10223} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10230};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10052} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9948} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10322};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10382} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10102} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10137};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10016 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9953} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10483};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3666} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9912};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9973} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10503} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10239};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10192} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9923} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10445};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10488} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10516} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10128};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10111} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9939} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10031};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[10]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10015} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10118};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10380} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10211} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10280};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10466} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10109} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10436};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9934};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10494} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10205};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9947} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10301} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10275};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[12]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10041} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10036} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9933};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10388} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10298} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10164};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9928} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10221};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10196} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10507} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10477};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10179};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10414} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10389} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10068};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10515);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10470} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10304} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10203};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10219} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10311} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10487};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10042} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10335} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10312};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9965} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9986} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10231};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10155} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10447} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10173};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10472 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10401} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9964} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10502};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10112} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10127} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9903};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10077} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10422} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10097};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10341} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10363} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9994};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10017} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10290};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10433 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10359} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10476} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10373};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9997} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10326} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10265};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10089} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10376} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10351};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9920} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10021} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10189};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10458 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10365} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10443};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10195} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10093} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10232};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10292} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10523} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9941};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3665);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10469} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10425} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10496};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10081} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10132} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10402};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10181 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[6]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10490);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10171} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10267};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10535} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10448};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10393} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10098} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10177};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10316} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10100} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9967};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10287 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22573);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10246} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10347};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9999} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10122};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3661);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10084};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[2]) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22567) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9981 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10336;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10354) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10266)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10134);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10481 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9989);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10480 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9919) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10404);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10254 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9906;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10314) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10188)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10043 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10449);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10079 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10468) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10327);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10367 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10022;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10464) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10110)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9978);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10157 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10212);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10379) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10344 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10056;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10446) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10035)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10534);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9916} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9976} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10242};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10303 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10187 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10532);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10034 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10009);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9952 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10166) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10438);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9972;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10255 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10051) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10123);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10385;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10143 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10119);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10169 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9957) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10440);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10252 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10519);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10020 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10261);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10092 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10510) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10357);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9938} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10185} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10209};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10106} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10460} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10491};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10374} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10129} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10032};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10138} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10410} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10529};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10063} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10162} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10331};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10473} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10096} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10361};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10399 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10299);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10434 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9983);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10115 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10018);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10151 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10397);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9911 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10161);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10296 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10269);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10408 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10536 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10227);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10358 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10073);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10202 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10257);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10395 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10451);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9969 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10121)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9988));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10525 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9944 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10427);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10215 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10083);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10200 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10346);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10424)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10289));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9987)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10479);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10539) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10387);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10207)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10076);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10486 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10204));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[32] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10372 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10146;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10497 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10345));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10243);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10377 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9996 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10492);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10355 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10463;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10277);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10437);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9977 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9918;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10467) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10533)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10302) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10352)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10222);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10145) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10144)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10010);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10249) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10117);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9936)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10420);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10241) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10108));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[32]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12770;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12051;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11490) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11386) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8144);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8231;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7993 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8521;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8481;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8322 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8573) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8247 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8107);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8591 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7854) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7877) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8054) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8344 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7972;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12416} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11613} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12556};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8539));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8348 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7761 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8095;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8385);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7829 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8303);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8038 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7781;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11650) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11457) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12044} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11233};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11353) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11257) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11891} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12799} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11686};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11254} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12751} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12489};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11894} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12571} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12634};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11420) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11323) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11520) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11501} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12446} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11647};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11961 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[5]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11222) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11218 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8327;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8364 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8560);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7864) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7678) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7940);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7903) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7739;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8325);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8479);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8436 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7805);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7701 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7860) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N771;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11712) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12309} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11803};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11379} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12156} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12607};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11506} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12280};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12363} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11657} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11370};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11752} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12453} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12516};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[37], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[36]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11785} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12749} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11858};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[37]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[37]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7951 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8688;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8187) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8610) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8358);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8753);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8319);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[18] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7898) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8428) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7911) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7691);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8367);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8788) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7755) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8512) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8652 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22714);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8284 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7736) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8683));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7950);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7992 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8053);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8141 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7910);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22705 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8608);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10213 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10082));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10364;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10400 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10520));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9954 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10493;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10465) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10325));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9943 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10426));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10167) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11925 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12149} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11492} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[36], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[35]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12260} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11470} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11532};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[36]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[36]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11383) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11287) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12834} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11755};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11617) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8039);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8643 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7764);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8091 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8020 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8740 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7994);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8267);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8152) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8401) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8351) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8778);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N770;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11781) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11487) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11677) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12083} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11418} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12229};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12589} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11729} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11512};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11995 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10459;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10008) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11255) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11744) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12341} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11844};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11454) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11350) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11550) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11536} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12484} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11680};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11269} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12100} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12821};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12722} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11762} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12284};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12401} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11160} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11932};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11646) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8355 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7975);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8650 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8565 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7683);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7946 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8276 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8700 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7843);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7918);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8082);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8422 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8558);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8762 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8527;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11855) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11416) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11320) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11963} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12871} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11826};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12756} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12620} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12650};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12849} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11351} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11870};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12526} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11289} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11542};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11407} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12668} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12184};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12547} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11280} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11568};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[31] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12869;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[30]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11317) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7974) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8217));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8460) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8594);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8684 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8165);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8556 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22699);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12471} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12626} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12059};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[35], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[34]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12427} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12866} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11441};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8540) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8292) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[17] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8204 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7717) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8072);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[17]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[35]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[35]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8300);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8522) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7776);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7743) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8477) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7998) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7857);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[16] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8328);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8639);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[16] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8092) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7858) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8579);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[16];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10023 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10524));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10403);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9917 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10313 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10174);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9979 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10175;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10065);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10006;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9925 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9985) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10475);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10285)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10152);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10293 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10158));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10381) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10105;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11708} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11185};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11819) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11516) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11709) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12119} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11460} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12262};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8625 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8242 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7798);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7871);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8490) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8729)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7968) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7709);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8299 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8069;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11921) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11615) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[1] & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10506;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22556;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11285) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11778) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11304} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12408} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12474};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12440} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11702} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11459};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12613} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11901} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12642};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7815) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7976 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8018) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7762);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8042);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7887);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8212 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12065} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12314} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12677};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11375) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12269} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11692} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11959};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[34], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[33]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12339} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12777} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11342};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[34]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[34]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[29]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[28] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12279;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11216) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11885) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11347) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12334} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12001};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11674) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12299} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12658};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11483) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11380) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11580) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11570} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12518} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11720};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12265} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11268} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12075};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12466} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11484} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12228};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10369 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10233));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10069;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10210 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10197));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10190 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10199;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10495) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10343);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10101 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9968));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10405) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9940) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11715 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11640} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11664} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11447) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12785} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11685} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11888};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8260) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8431);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8078);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8746 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8308);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8132);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7719 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8697) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8614)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8667) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8372);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8001 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8235);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7862) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7891;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7670) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8607);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7778 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8034 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7896 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8123);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8439);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8708 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7851;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11988) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12376) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11881;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11450) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11548) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12151} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11188} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11920};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12107} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12035} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11306};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12291} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12791} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12043};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12256} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11235} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11261};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11282) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12407} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11945} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11310};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11511) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8380 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7797) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7708 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8601);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8090) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7966 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8782) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8102);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8681 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44095);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11851) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7789);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7806 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8386 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8630);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8432 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8576) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8249);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8229) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8613)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8518) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8714 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8056 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8309);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8538 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8772);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8147 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8495 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7878;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12055) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11741) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11638} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11493} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12300};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12082} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11880} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12619};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12765} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11843} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12588};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12683 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[27]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[26] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12830;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12836) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12011} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11172} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12491};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12435} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11499} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11417};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11833} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11319} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12581};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[33], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[32]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12460} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12691} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11476};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7763);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8083;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8044) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8252 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8010);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8293);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8258 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7971);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8234);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[15] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8112) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8545) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8151);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[15]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[33]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[33]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8314 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8784);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8468) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7726) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7682);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8420);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[14] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7945 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8507) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7793));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10450 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10317));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10000) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10457;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10178 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10044));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10216) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10120;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10412 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10273 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10333) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10194);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43743) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43757)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10156) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11620);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11513) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11412) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11611) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11606} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12552} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11757};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11706) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11918) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12021) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12825} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12687} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12072};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11890} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12837} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12657};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11952) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11644) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11814) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12411) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8458 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8209);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7938);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7978);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8715 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8596);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8559 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8169);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7784) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8754 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8520;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12120) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11956} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11919} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11262};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11339} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12441} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12118};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12798} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11854} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11649};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11812} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11612};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11345) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12034} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12729} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12660};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8062);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8286) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8188 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8172);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7732) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7820) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7894 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8160) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8706);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8655 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12086) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7863 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7811);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7676) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8541) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7957) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7816);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8636 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8394;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12181) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12186} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11672} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12614};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11480) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11373;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11228} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12549};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11777) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11882) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11671) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11529} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12333} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11371};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12367} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12150} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12870};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11679} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12627} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12448};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12596} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12415} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11427};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11181) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12561} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12168} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12122};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11574) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12831} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11772} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12758};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12192} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11449} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11194};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[32], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[31]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12094} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11602} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12813};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[32]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[14]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[32]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11637) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11409) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12481} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12306} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12383};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12593 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[25]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[24] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43395;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12741) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11477) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12202} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11924};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8771 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8537);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8713);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8598 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8430 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8003);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8246);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7703);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8055 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8323) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8012);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8143 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44079);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11721} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12483} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11500};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11654} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11466} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12236};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11248) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11621} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11393} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11723};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11584} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12351} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11388};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11802} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12530} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11549};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[31], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[30]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12221} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11967} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11224};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8280) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8379) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7752);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8624);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8340 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8770);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8086 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8006);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7921 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8185) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[13] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7965);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[13]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[31]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[31]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8640 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8118));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8356);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8483 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8466);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8071) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8027) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7771) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8469);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[26] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8218 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8701);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[26]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8088) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8362) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7696 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8124) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7970);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7848);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8738);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8426)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7735);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[25] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7799) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8139)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7873) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8243);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[25]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12786) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8647) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7835);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8339 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7890);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8109);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8334) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7672) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8302);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8658 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8410);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[24] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8036 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7779);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[24]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[41] = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[42];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8400) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7786);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8227) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8127) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8474;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8767 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7855) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7953 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7698);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[23] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8190);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12817) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12850) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[41], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[40]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11730};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[23]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[41]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[41]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7814) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8396);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8543);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8255);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8125 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[22] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7886) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8210) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7919);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11196) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12270;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11423) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11165) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12760));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11263) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11771} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12695};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[40], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[39]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11886} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11352} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12479};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[22]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[40]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[40]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8207 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8698) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7839);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8175);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8711) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8664) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[21] = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8629 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8101) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7819) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8523;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[39], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[38]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11953} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12116} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12684};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[39]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[39]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8501 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8128 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8376;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7962);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8725) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8587);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8065 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8447);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7750) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8622) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[20] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8779);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[38]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[38]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11700) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9907 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10394));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10183) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43770;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10256 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10124));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43769 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43761;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43747) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43739) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11523 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11545) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11848) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11410;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11957} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12582} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12609};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11984) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11641) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12146) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7989 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7767);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8310 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8561);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8756 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7679 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7838);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8418 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7942);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8504 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8148);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8075 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8213);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8174);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7790 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8045;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12246) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11298} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11793} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12254};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12475} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12403} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12185};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11739) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11950) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12052) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12862} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12717} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12108};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11187} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11756} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12519};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12663} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12274};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11916) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12117) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12212) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12648} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11710} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11563};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22572 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12412);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12040));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11607) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11874} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12224};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11810) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7748 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7901);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8375 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8485);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8099 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8620 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8004);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8134);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7706);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8446 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8679);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8064 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7817;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12310) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12020) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11871} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12508};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12437} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11453} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12223};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11994} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11962} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11535};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11275} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11687} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12053};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12423} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11434};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8251) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7883);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7718);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8304) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8461)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7753) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7775) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8206);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8167) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7782)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8275);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11313) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11239} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12386} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11344};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12388} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12115} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11395};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12803) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11543) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11770) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11531} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11161} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11718};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11201} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12170} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11977};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11360} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12162} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12136};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[30], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[29]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12555} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12318} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11577};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7693);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8011) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7935) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7727 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8345) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7824) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8161;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[12] = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8033) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7705) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8656;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[12]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[30]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[30]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11795} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12029} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12551};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11878) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12469;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11993} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12669};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11703) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11982) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8298 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8265 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8028);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8470 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8703);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8405);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7892);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7983 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8084 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8546);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7826) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8119) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7932) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8158);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7684 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8568;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12370) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11773) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11485} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11180} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12752};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11411} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11704} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12257};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11643));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11667) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12177) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12277) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11333} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11837} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12292};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12068} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11488} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12788};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12004} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11227} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11569};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12692} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12308} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11725};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8094 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7982);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7769));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8383;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8581);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8717 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8232) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7788) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8315);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8329 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8437) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8058)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7787) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8416);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11372) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11619} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12455} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12690};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12505 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[23]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22582;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12655) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12865) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12344} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12775} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12525};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12018} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12209} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11207};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9990 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10482));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10235) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10229;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10337 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10201));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10452;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10099) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9966));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12350;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11314} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12089};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11603) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11842) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12868} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11472} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11337};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12736} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11987} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11780};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11174} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12703} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11948};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[29], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[28]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11168} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12857} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11939};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8443);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7738) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8324) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8478) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8365);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7856));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8163);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[11] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7695 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8189) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8673));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[11]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[29]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[29]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11212) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12707) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11665) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11969} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12155} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12515};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8616 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8154);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8642);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8503);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8509) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7766) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8488);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8019);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[8] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7924 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7723) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8602) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8113);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11947) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12144) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11743;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11748} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12723};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12084) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11734) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11846) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7960);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8342);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7744);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8177 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8427 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7939) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8052) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8283;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8338 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7754);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8535 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7801 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8732 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7874);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8590 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7711);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8454 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8198;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12432) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12402} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11451} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12819};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12143} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12705} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11525};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11836} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11264} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12584};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12340} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12725} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11346};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11443) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12493} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12592} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12338};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12245} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11249} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11821};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20]) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[20] ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11979;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12562) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12244) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12337) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12050) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11910} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12679} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12542};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12506} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12822} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11873};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12399) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12210) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12307) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11362} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11521} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12323};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11265);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11912) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12674} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11329} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12030};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12017) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11806) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12113) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12789} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11217} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12179};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12740} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11782} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12538};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11328} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12293} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12616};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12038} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11605} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12759};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10071 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9931));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18] = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N9962) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10047;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18] & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12138} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12859} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12352};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12173) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12617);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12275) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12319} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11786} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12711};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11940);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11742) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12494) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12366) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11980) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12080) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11634} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11949} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12573};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12467} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11823} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12568};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12459) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11875) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12258);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11943) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12701} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11552} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12066};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12438} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12858} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12604};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12389} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11396} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11591};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12327} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11558} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11913};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11301} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11642} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12076};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12375} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11805};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11387} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11765} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12527};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11909) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11508} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12807} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12686};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12566} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12024} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11589};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12710} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12536} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11747};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[28], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[27]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11740} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12502};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8226);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8208) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7884) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8228 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8200);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8557 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8498);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[10] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7673) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8686) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[28]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[28]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12771) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11278) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11731) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11763} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11576} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12148};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11507) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8171 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8769);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7728) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7700 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8589);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8421);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7925) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7913) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8262) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8081);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8316);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7833 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8133) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8237)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8550) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7844);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11850} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11960} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12124};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12281} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11283} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11859};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12622) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11571) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11382} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12731} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11566};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11976) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12832) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8615) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8742) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7821) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8731);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8606)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8381) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8452);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[6] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8552 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8068) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7930) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8787);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11341) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12797} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11193} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11378};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12329} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11544} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12315};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12601} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12061} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11626};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12745} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12357} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11788};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[27], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[26]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11556} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12511} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12326};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8079 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8553;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8253 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8651) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8442) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8273) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7899) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8129);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7999) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7861) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[9] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8330));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[9]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[27]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[27]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11804) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10417 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10279));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10148) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10013) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10258;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10315) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10390) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N10176);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11978);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11713) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12524) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11270));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12046) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12141) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11256} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12503} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12216};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12429) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12240) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12335) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11402} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11557} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12358};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11628} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12398} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11436};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12172} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12360} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11176};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12653} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11335};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12468) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12410} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12794} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12200};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11754} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12158} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12558};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11322} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12842} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11896};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12042) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12681) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11635) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11421} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12382} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11184};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8272);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8564) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8361);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8577 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7734) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8555;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7772 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7991);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[5] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7690 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7852) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8709) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11405) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11179) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12721} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12078} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12557};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11579} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11955} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12346};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12637} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12096} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11659};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12395} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12779} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11827};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[26], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[25]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11363} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12142};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8445 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8722);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8678);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8063) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8153) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8649 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8021);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7765 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8741);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8236 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8195) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8043;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[8] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7888) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8291) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8402) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[8]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[26]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[26]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7740);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8026) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8510);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8002 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8532 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8567 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8269) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8566);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8180 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7729) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7794;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[7] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8277 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7955) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8763);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11872) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12396) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12015) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12110) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11666} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11985} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12611};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11489);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12737} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11775};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11876);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12207) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12531} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12253} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11828};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12433} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11445} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12247};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11211} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12211} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11404};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11364} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12595};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11675} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12111} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12443};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12106) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11847} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11561};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11163} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11354} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11934};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12532) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12739) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11697) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12009} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11811} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12548};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12492) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12304) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12272) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12077) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11868} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11442} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11292};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12746} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11173} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11258};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11251} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12026} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12218};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11989} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12182} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11853};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12682} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12145} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11716};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8575 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8216);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8089 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8140) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8593) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7757);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8735 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7849) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7715);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8349 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7900) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8197 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8146) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8374);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7915 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8388);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22659 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8494);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22587) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11474) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11303} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12829} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12374};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12194} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12591} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11616};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12670} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11695};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12430} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12815} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43997};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[25], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[24]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11401} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12574} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12178};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[25]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[7]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[25]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8611 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8205);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7876 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8648) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8282);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8166);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7952);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7947) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8730) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7710);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7872 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8009);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8453) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7792) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8104) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8785);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[6] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8070 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22592) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11941) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11245) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12169) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12191} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12714} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11178};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11197} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11971} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12384};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12801) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11691));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12361) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12456) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12019);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11681) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12550) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11590} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12394} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12537};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12033} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12062} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12782};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11220} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12748} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12800};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12712} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11182} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11750};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11429} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11614} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12864};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8768);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8363) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8097)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8467) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7885);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7830) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7803) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8661) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8312);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7783) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7777) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8519) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8584);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11767) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11539) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12183} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12297} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12000};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11463} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11884} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12623};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12010) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11311) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11801} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12365} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12477};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12231} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11652} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11236};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11391} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12697} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12164};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12851} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12462} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43976};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[24], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43957} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43935} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43964};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[24]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[24]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11318));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12652) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12238) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12425) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12733} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11863} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12025};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12171) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12520) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12332) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12139) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12780} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11208} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12643};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12252} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11840} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12586};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12754} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11830} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12578};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11998} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11790} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12545};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12863) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12764} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11234};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12235) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11839) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8023 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8008);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7677) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8514) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8582);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8462) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8150);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8233) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8480);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8440) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7810);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7958 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11526} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11791} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11601};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12539} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12659};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12074) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11369) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11419} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11992} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12512};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11495} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11682} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12267};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12014} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12418} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11430};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12497} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11732} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11169};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43982} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43938} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43944};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8397 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8145;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8110 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7865 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7917);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8360) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7760 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44116);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8050) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8263) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8666) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7990);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8301 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7882);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43970) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43954) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8215) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43941);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43985} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43987} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43994};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14822 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14841);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12393) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12487) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11276) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12575) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11210));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11627} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12431} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12567};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12470);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12302) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12773} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12013} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11479};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11425} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12196} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11456};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12612} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11636} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11610};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12081} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11800} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11599};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11505) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12201) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12406} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12371} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11215};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12667));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12704) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11206) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12414} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12719} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12587};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7926 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8644);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8692) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8696)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8415 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8285 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8294);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8743) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8403) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8164 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8076) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8562) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7979) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11905) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11662) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11408} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12507} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11225};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12336} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11538} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11340};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12767) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12313);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12268) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12454) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11237} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11904} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12060};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12104));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12205) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12535} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12761};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12226} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11199} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11231};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12405} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11305} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12379};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11274) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12554} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12045} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12230};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12356) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8502 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8721);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8638 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8176);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8702 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7967) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8765) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8183);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8781 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8716 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7800) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8392) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8724) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8473) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8278 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7846);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8111 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8529);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8335)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7685) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7749);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12166)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11972) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11727) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12750} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11746} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12580};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11784} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11758} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12522};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12482) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12264) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11175) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12424) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12517) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12606) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11660} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12461} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12602};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12090) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12809) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12546) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12747));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12359) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11705);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12328) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12808} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12232} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11514};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11247} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11917};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12656} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12167} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11171};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11809} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11555} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12559};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11528} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12321} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11582};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11400) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11267} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12700} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11458};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12570} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12744} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12161};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11540) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12828) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11776 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11415} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11648} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12706};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12421) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11930);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12301} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11973} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12008};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11338) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11385} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12188} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11845};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11397} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11572} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12343};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12872} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12125} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11929};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12838} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11892} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12091};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11307} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11502} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12276};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12135) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11440) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12757} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11592} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11564};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12486} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11530} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12303};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12298) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12176} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12688} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11722};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22586) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11799) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12039) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11567) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12400} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12220} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12036};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11376} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11349} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12153};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12311} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12121} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11316};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12085} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12802} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11277};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[19], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11856} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12056} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12597};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8106 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7687);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8350 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8408);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7908);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8645) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8352) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8450 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8025) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8224) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8694);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8547) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7804)) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7770) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7680);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8506) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8524;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[1] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7943) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7897) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7937);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11272} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12449} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11468};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12768} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12047} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12239};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[20], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[19]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11242} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12563};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[19]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8627 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8192);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7812 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7694);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7841 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7859);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8059) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8526) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8719) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8737);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7692) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7813) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7870);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8067;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7780) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8115)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8399) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7831);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[2] = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8395) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8542) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7920);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12732} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11774} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12204};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[21], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[20]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12533} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11203} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11551};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[20]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8239 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8617);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7987);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8391 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8434);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7675) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8331) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8413) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8040 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8035);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7742 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7995);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8317) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7785) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8755) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[3] = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8157 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8126) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8626) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8612;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[21]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43947} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43960} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43990};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[21]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14601 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7697 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7931) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8393) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8230);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8250 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8041);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734 = ((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7916 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7725) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8764) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8747;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8037) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8307)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7934) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8734);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8727 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43963) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43949);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43993} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43967} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43973};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14522 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12103) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11633) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11867) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11639} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12028} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11834};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11191} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11166} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11966};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12325) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12540) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12728} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12213} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12392};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11471) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12165) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12793} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12348} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11632};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11241) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12874);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12485) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11330);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12572) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11462} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12097} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11284};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12772} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11527} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12296};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12509} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11946};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11331} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12621} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12243};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11737} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12499} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11768};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11937} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12693} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12673};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12846} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12665} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11900};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[18], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12629} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12810} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11655};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8429 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8528;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8569) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7949) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8223) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7902) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8354) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8048);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8669) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8777) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8486) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8531);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8105 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7802 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8135);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8371) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8633)) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7845) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8621);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[0] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8586 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N8016) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7961));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[0]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14673 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11694) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11936) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22590) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12387) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11448} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11260} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11825};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11308) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12543) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12843} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12444} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11696};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12390) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12852} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11954} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12420};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12523);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11820} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11302} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11749};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12445} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12263} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12676};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11464);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12734) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12600) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11392));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12022} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12105} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11357};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11519} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12529} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12288};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11728} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12496} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11698};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11688} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12639} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12458};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11764) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12007) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22593) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12447) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12784} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12615} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11439};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12233) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22579) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11534) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12123);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12638) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12635) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12576));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12450) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12513) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12320);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12603) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11676} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12128} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11321};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12498} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12636} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12599};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12685} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11433} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12709};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12565} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12079} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11281};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12442} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11253} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11465};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12824} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11877} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12134};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11547} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11295} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12316};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11509} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12464} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12283};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11560} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12331} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11986};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11437) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11719} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12206} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11494};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22577;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11658) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12353) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22574 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11944);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12569) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11164} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12651} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11733};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12159);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11481) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12664) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11413));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12630) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11553 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11170 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22561);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11293) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12689) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11668));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3662} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12860} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12696};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11914} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11355} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12428};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12671} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12867} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11991};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11533} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12242} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12305};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12095} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11624} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11336};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12250} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12480} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11673};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12796} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11588} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12355};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12472} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11491} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12016};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11594) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11761) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11365) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12294) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11879} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12073} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12608};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12514) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11835) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43396;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44110;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12070) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12354);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11915) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12510) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12295));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12436} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12255} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12776};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12234} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11707} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11238};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12854} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12618} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11906};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12647} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11645} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11670};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12071} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11325} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12099};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11970) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12198) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11663} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11486} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12114};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11503) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12769) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12419) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11432));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11724) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11861} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12826} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11299};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11498} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12271} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11983};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11902) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22585) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12133) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12064} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11869} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11205};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11849} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11361} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12594};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11618} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12140} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12385};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12259} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12735} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11266};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15031 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12208} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11923} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12848};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11794) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22588) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12261) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12649} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11309} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11290};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11377);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12720));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11565) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11209} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11244} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12473};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12391} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11399} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12833};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12708} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11273} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11745};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12037) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12426) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11864) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11630) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11622);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11177) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12322) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12478));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12109} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12290} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12641};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12820} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12023} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12088};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11887} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12175} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12625};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12102) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11690) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11593} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11435} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11711};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12465} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12662} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12716};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12806} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12743} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11783};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14853;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11999);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12058} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12422} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11938};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11933) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12713) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12163) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12101} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11438} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11911};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11753} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11684} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12452};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12451) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12227) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12804));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11760) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22578) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12003) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11332} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11701} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11522};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12364} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12214} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11367};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22581) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12067) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12628} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12702};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11899) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11990) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12129) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12362));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12324} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12490} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12504};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12841} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12856} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11895};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11600);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12534 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11223));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11829) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12137} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11653} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12680};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12632} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12778} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11824};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11965) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12579);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11631 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12219);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[1]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12835} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[19]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3], DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11889} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11343};
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11288 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11183);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[1] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12488) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12032) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N12839));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[1] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N11504 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[3] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14697 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15072) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14944);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14690) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14733)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14615);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15041 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14745) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14625);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[5] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[6] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14871 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14679) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14572) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14623)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15069);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[7] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14529 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14924) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14797);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[8] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14807) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14604)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15055);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[9] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[10] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14724 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14530) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14974);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14940;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15016 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14887) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14763);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[11] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14777) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14751)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14658);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[12] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[13] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14904 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14707) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14582;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14565 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14627) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15075);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[14] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[15] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14834 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14638) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15083);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15057) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14534)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[16] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14965 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14882) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14756);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14635;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[17] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14621 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14992) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14867);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14599 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14718 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14845);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14918 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14545) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14792);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14970 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14650 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14772);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14847 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15048) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14719);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14895 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14577 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14699);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14773 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14971) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14634 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14861;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14823 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14948);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15074 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14628);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14749 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14874);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14998 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14554);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14682 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14801);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14927 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14607 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14728);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14855 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14978);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14535 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14661);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14909 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14779);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14586 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15034);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14710 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14836);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15087 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14956);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14758 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14931)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14812));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15011 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14885);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14692 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14562);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14934 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14813);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14616 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15066);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14646)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14515));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14865 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14736);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14987 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14541);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14671 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14788);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14914 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15043);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14923)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14795));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15052)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14922);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14558) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15001);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14700 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14712) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14694)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14566);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837 = !((N22531 & N22593) | N22648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14596 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14716);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14966 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14843);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15006 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837) & (!N22536)) | N22534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43813;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14706 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14543 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14738;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14990 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14985 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14580;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[48] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837 & N23056) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837) & N21801));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[48] & N21766);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22752);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219 | N19980);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14787 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14849);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14794;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14783 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14722 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14774) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808 = !(((!N22564) & (!N22562)) | (!N22566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[28] = N22489 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[28] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14556 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14999));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14826 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14875;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14703 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14594) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14750;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[29] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808 & N22387) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14808) & N22385);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[29] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14589 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14938;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15038 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14620 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14896 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14761 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14911);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14951 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15028;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14644 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14579 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14631) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771 = ((!N22566) & (!N22571)) | (!N22569);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908 = !((N22504 & N22644) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14771);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[40] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908 & N22402) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908) & N22404));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[40]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14693 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14563));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15012;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14858 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14886);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14714) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14832)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14958 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14600;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14840 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14846 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14817;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[41] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908 & N22409) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908) & N22411));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[41]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14617 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15067));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14760 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14643 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14688) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14767);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14725);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14872);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43441 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15015 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14590);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15020 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14967;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14893) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14945)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14821);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426 = !N22510;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14746) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14799)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14680);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14605) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14660)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14531);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15039 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15033) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15084)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14645) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14622)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14888 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14878) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14752);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433 = ((!N22512) & (!N22583)) | (!N22581);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43426 & N23029) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43433);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[43] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585 & N22366) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585) & N22368));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[43]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14881 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14935 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14814));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[42] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585 ^ N22319;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[42]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14669 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[46] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837 ^ N22392;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[46] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15045 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14915));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14739 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14789;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14619 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15040) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14672;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[47] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837 & N22439) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14837) & N22437);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[47] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14564 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14555;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15014 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14803 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[44] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585 & N22453) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585) & N22451);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[44]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14866;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14869);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14737 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14588);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14542 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14988));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43432 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14994) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14689)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43449);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43446 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43424 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43438;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14585;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434 & N22330) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43434) & N22332));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43448);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14759 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14641));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14782 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14665 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14903) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[39] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908 & N22395) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908) & N22397));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[39]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14528 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15088 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14957));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[38] = N22361 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14908;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[38] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14838 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14711));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14557 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14975)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14980 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14982;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14859 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14667 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14963;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14602);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15025 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14649 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14666 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15089);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14775;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14830 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14902;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14537 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14526 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15050) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14972);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14959 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14900 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14950) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14827);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521 = ((!N22520) & (!N22600)) | (!N22598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662 = !((N22558 & N22646) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14521);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662 & N22482) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662) & N22484));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[37] = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44122;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[37]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14587 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15036));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15010 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14609 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14753;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15061 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15003 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14883;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[36] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662 & N22344) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662) & N22342);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[36]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14910 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14780));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43800 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43804 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14550;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662 & N22351) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662) & N22349);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43808);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43811 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14663 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14536));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817 = N22373 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14662;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43817);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14571 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063 = !(((!N22526) & (!N22524)) | (!N22528));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[32] = N22416 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[32] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14979 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14856));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15000 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14729;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14877 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14943) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14608;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[33] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063 & N22432) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15063) & N22430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[33] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15059 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14928));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14630 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15079 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14768) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929 = !(((!N22510) & (!N22508)) | (!N22512));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[31] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929 & N22358) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929) & N22356);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[31] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14964 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14802 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14683));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[30] = N22378 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14929;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[30] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14701 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14578));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14652 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15023) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14525 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14897) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14810;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732 = !N22531;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[25] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732 & N22442) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22732) & N22444));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[25]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14614 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687 = !(((!N22518) & (!N22516)) | (!N22520));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[26] = (!N22304) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[26]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14629 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15076));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15024 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14949) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14899 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14824) ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14986;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[27] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687 & N22421) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N14687) & N22423));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2] = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22595 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[27]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15920)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15959);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15945);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15967) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15987);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15978)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15917);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8] | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15994) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15923);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12] | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15931) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15950);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15941) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15972);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15962 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15913);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16] | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15960) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15980);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15970 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15989) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15983);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15911) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15937);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15949;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0] = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43335;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43365);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43353 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43361);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15954;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15982 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15934) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15928);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15984 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15963));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15921;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15938 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15992) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15958);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43367) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43337);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15946 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15944));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15976) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15956 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43345);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43706) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43715);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[1] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43346));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15990;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15926;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15996) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43708)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43717);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43693 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15953));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952) & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43689)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43696);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N43713;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[22]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16087) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16139));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N541;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15969 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15935));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072 = (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N44129) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16062);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4] = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16072) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15952) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16063));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16107) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16144 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N542 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N543);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[0] | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16065);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3] = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16069 ^ DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16170));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670 = (N23330 & N20260) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N701);
assign x[22] = (N23314 & N23328) | (N23321 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[3]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[5]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[1]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[0]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[19]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[21]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[15]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[17]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16108));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16229) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[11]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[13]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[7]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[9]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16113 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16133));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584 = (N23335 & N20547) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N700);
assign x[21] = (N23316 & N23328) | (N23323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16100) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16188));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16241 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16176) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16109));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16197) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16126));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16195) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16214) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16147));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16169));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16234 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16099));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668 = (N23331 & N20392) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N699);
assign x[20] = (N23319 & N23328) | (N23326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16222) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16154));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16140) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16231));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16163) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16093));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16196));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16161) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16203) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16132));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16201 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16221));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667 = (N23332 & N20454) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N698);
assign x[19] = (N23318 & N23328) | (N23325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16240 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16182) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16162));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16124) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16220) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22599) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16202));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16166 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16189));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666 = (N23333 & N20350) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N697);
assign x[18] = (N23314 & N23328) | (N23321 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16175 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22600);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16146) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16104) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16125));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16091) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16187) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16168));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16130 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16155));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665 = (N23336 & N20537) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N696);
assign x[17] = (N23315 & N23328) | (N23322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16105 | (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22596));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16114) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16092));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16212) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16153) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16131));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16096 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16120));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664 = (N23330 & N20444) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N695);
assign x[16] = (N23318 & N23328) | (N23325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16235) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22597) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16213));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16181 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16119) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N22598) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16098));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16218 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16207));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663 = (N23335 & N20557) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N694);
assign x[15] = (N23317 & N23328) | (N23324 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16186 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16138));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662 = (N23331 & N20414) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N693);
assign x[14] = (N23317 & N23328) | (N23324 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16151 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16228));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661 = (N23333 & N20360) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N692);
assign x[13] = (N23314 & N23328) | (N23321 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16118 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16159));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660 = (N23335 & N20434) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N691);
assign x[12] = (N23319 & N23328) | (N23326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16206 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16090));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659 = (N23333 & N20481) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N690);
assign x[11] = (N23319 & N23328) | (N23326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16136 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16180));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658 = (N23334 & N20471) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N689);
assign x[10] = (N23316 & N23328) | (N23323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16225 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16111));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657 = (N23334 & N20424) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N688);
assign x[9] = (N23315 & N23328) | (N23322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16158 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16219);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16200));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656 = (N23333 & N20587) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N687);
assign x[8] = (N23319 & N23328) | (N23326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16129 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655 = (N23332 & N20577) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N686);
assign x[7] = (N23314 & N23328) | (N23321 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16216 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654 = (N23334 & N20370) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N685);
assign x[6] = (N23317 & N23328) | (N23324 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16150 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653 = (N23332 & N20491) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N684);
assign x[5] = (N23316 & N23328) | (N23323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16239);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652 = (N23330 & N20567) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N683);
assign x[4] = (N23317 & N23328) | (N23324 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16172 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651 = (N23330 & N20501) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N682);
assign x[3] = (N23315 & N23328) | (N23322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650 = (N23334 & N20597) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N681);
assign x[2] = (N23316 & N23328) | (N23323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16192);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649 = (N23332 & N20607) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N680);
assign x[1] = (N23318 & N23328) | (N23325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16121 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648 = (N23331 & N20617) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N679);
assign x[0] = (N23318 & N23328) | (N23325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487 & (!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647 = a_exp[7] & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N639;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[30] = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N759 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N580) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16646 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N647);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468 = !((N23333 & N21461) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__219 & (!N23330));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16468 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426);
assign x[29] = (N23319 & N20199) | (N23326 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422 = !((N23332 & N21468) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16422 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426);
assign x[28] = (N23314 & N20199) | (N23321 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675 = !DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482 = !((N23335 & N21042) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N675));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16482);
assign x[27] = (N23318 & N20199) | (N23325 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436 = !((N23335 & N21116) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[3]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16436);
assign x[26] = (N23315 & N20199) | (N23322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391 = !((N23331 & N21231) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__215[2]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16391);
assign x[25] = (N23315 & N20199) | (N23322 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449 = !((N23331 & N21208) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16178));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16449);
assign x[24] = (N23316 & N20199) | (N23323 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405 = !((N23334 & N21450) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16452 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16142));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16405 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16426);
assign x[23] = (N23317 & N20199) | (N23324 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540 = (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N661 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N654) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N666;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N657 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N664 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N668);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16578 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16560);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16540 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16547);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N653 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N651) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N658);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N660 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N659) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N667);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16570 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16542);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530 = ((N20988 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N645) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N646) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N640;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N641 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N642) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16530);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N643 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N644);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16565 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16557 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N648) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N655);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N663 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N656);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16576 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N649 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N650) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N652);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N665 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N3584);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16556 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16572);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563 = DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16535 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16558;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16575 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16563);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7373 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7196);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757 = !(DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7297 | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N7131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577 = !((DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757 & a_sign) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N757) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N15829));
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16612 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N577) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N487) | DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__82);
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607 = (!N20253) | (DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16545 & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16532);
assign x[31] = !((N23336 & N19976) | ((!N23336) & DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_N16607));
reg x_reg_30__I4228_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I4228_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[30];
	end
assign x[30] = x_reg_30__I4228_QOUT;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[0] = x[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[1] = x[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[2] = x[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[3] = x[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[4] = x[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[5] = x[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[6] = x[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[7] = x[7];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[8] = x[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[9] = x[9];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[10] = x[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[11] = x[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[12] = x[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[13] = x[13];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[14] = x[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[15] = x[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[16] = x[16];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[17] = x[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[18] = x[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[19] = x[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[20] = x[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[21] = x[21];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[22] = x[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[23] = x[23];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[24] = x[24];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[25] = x[25];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[26] = x[26];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[27] = x[27];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[28] = x[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[29] = x[29];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[31] = x[31];
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__42[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__195[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__197[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__201[49] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_0_inst_inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urTzQg/eohpI : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



