/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:24:20 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module cynw_cm_float_cos_inst_cellmath__231_0_bdw1114505291_bdw (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__21,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire  inst_cellmath__46;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__66,
	inst_cellmath__67,
	inst_cellmath__68,
	inst_cellmath__69,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__200,
	inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire  inst_cellmath__219;
wire N491,N492,N493,N494,N548,N549,N550 
	,N551,N552,N583,N585,N594,N595,N597,N598 
	,N599,N600,N601,N602,N603,N604,N605,N606 
	,N607,N608,N609,N610,N611,N612,N613,N614 
	,N615,N616,N617,N618,N619,N620,N621,N622 
	,N623,N624,N625,N626,N627,N628,N629,N630 
	,N631,N632,N633,N634,N635,N636,N637,N638 
	,N639,N640,N641,N642,N643,N644,N645,N646 
	,N647,N648,N649,N650,N651,N652,N653,N654 
	,N655,N656,N657,N658,N659,N661,N662,N663 
	,N664,N665,N666,N667,N668,N669,N670,N671 
	,N672,N673,N674,N675,N676,N677,N678,N679 
	,N680,N681,N682,N683,N684,N685,N686,N687 
	,N688,N689,N690,N691,N692,N693,N694,N695 
	,N696,N697,N698,N699,N700,N701,N702,N703 
	,N704,N705,N706,N707,N708,N709,N710,N711 
	,N712,N713,N714,N715,N716,N717,N718,N719 
	,N720,N721,N722,N723,N724,N725,N726,N727 
	,N728,N729,N730,N731,N732,N733,N734,N735 
	,N736,N737,N738,N739,N741,N742,N743,N744 
	,N745,N746,N747,N748,N749,N750,N751,N752 
	,N753,N754,N755,N756,N757,N758,N759,N760 
	,N761,N762,N763,N764;
cynw_cm_float_cos_inst_blk01_cellmath__39_bdw1114505291_bdw cynw_cm_float_cos_I0 (.inst_blk01_cellmath__39_out0({N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597}), .inst_blk01_cellmath__39_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_cos_inst_cellmath__42_0_bdw1114505291_bdw cynw_cm_float_cos_I1 (.inst_cellmath__42_0_out0({inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6], inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__42_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__48_bdw1114505291_bdw cynw_cm_float_cos_I2 (.inst_cellmath__48_out0({N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684}), .inst_cellmath__48_in0({inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__48_in1({N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623}));
cynw_cm_float_cos_inst_cellmath__58__24__bdw1114505291_bdw cynw_cm_float_cos_I3 (.inst_cellmath__58__24__out0({N493, N492}), .inst_cellmath__58__24__in0({N708, N707}));
cynw_cm_float_cos_inst_cellmath__61_0_bdw1114505291_bdw cynw_cm_float_cos_I4 (.inst_cellmath__61_0_out0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17], inst_cellmath__61[16], inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__61_0_in0({N492}), .inst_cellmath__61_0_in1({N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684}));
INVXL cynw_cm_float_cos_I5 (.Y(inst_cellmath__115__W1[0]), .A(inst_cellmath__61[16]));
cynw_cm_float_cos_inst_cellmath__195__80__2WWMM_2WWMM_bdw1114505291_bdw cynw_cm_float_cos_I6 (.inst_cellmath__195__80__2WWMM_2WWMM_out0({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0], inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0], N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742}), .inst_cellmath__195__80__2WWMM_2WWMM_in0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17]}));
cynw_cm_float_cos_inst_cellmath__198_0_bdw1114505291_bdw cynw_cm_float_cos_I7 (.inst_cellmath__198_0_out0({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17], inst_cellmath__198[16], inst_cellmath__198[15], inst_cellmath__198[14], inst_cellmath__198[13], inst_cellmath__198[12], inst_cellmath__198[11], inst_cellmath__198[10], inst_cellmath__198[9], inst_cellmath__198[8], inst_cellmath__198[7], inst_cellmath__198[6], inst_cellmath__198[5], inst_cellmath__198[4], inst_cellmath__198[3], inst_cellmath__198[2], inst_cellmath__198[1], inst_cellmath__198[0]}), .inst_cellmath__198_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__198_0_in1({inst_cellmath__115__W1[0]}));
cynw_cm_float_cos_inst_cellmath__203_0_bdw1114505291_bdw cynw_cm_float_cos_I8 (.inst_cellmath__203_0_out0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__203_0_out1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__203_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__203_0_in1({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17]}), .inst_cellmath__203_0_in2({inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0]}), .inst_cellmath__203_0_in3({N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742}), .inst_cellmath__203_0_in4({inst_cellmath__115__W1[0]}));
cynw_cm_float_cos_inst_cellmath__201_0_bdw1114505291_bdw cynw_cm_float_cos_I9 (.inst_cellmath__201_0_out0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}), .inst_cellmath__201_0_in0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__201_0_in1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__201_0_in2({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0]}));
cynw_cm_float_cos_inst_cellmath__200_0_bdw1114505291_bdw cynw_cm_float_cos_I10 (.inst_cellmath__200_0_out0({inst_cellmath__200[48], inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0], inst_cellmath__200[24], inst_cellmath__200[23], inst_cellmath__200[22], inst_cellmath__200[21], inst_cellmath__200[20], inst_cellmath__200[19], inst_cellmath__200[18], inst_cellmath__200[17], inst_cellmath__200[16], inst_cellmath__200[15], inst_cellmath__200[14], inst_cellmath__200[13], inst_cellmath__200[12], inst_cellmath__200[11], inst_cellmath__200[10], inst_cellmath__200[9], inst_cellmath__200[8], inst_cellmath__200[7], inst_cellmath__200[6], inst_cellmath__200[5], inst_cellmath__200[4], inst_cellmath__200[3], inst_cellmath__200[2], inst_cellmath__200[1], inst_cellmath__200[0]}), .inst_cellmath__200_0_in0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}));
cynw_cm_float_cos_inst_cellmath__17_0_bdw1114505291_bdw cynw_cm_float_cos_I11 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__46__15__bdw1114505291_bdw cynw_cm_float_cos_I12 (.inst_cellmath__46__15__out0({N491}), .inst_cellmath__46__15__in0({inst_cellmath__42[7], inst_cellmath__42[6]}));
cynw_cm_float_cos_inst_cellmath__46_0_bdw1114505291_bdw cynw_cm_float_cos_I13 (.inst_cellmath__46_0_out0(inst_cellmath__46), .inst_cellmath__46_0_in0({N491}), .inst_cellmath__46_0_in1({inst_cellmath__42[8]}));
cynw_cm_float_cos_inst_cellmath__21_0_bdw1114505291_bdw cynw_cm_float_cos_I14 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__83__62__bdw1114505291_bdw cynw_cm_float_cos_I15 (.inst_cellmath__83__62__out0({N494}), .inst_cellmath__83__62__in0(inst_cellmath__46), .inst_cellmath__83__62__in1(inst_cellmath__21), .inst_cellmath__83__62__in2(inst_cellmath__17));
cynw_cm_float_cos_inst_cellmath__19_0_bdw1114505291_bdw cynw_cm_float_cos_I16 (.inst_cellmath__19_0_out0(inst_cellmath__19), .inst_cellmath__19_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_cos_inst_cellmath__24_0_bdw1114505291_bdw cynw_cm_float_cos_I17 (.inst_cellmath__24_0_out0(inst_cellmath__24), .inst_cellmath__24_0_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_cos_inst_cellmath__69_0_bdw1114505291_bdw cynw_cm_float_cos_I18 (.inst_cellmath__69_0_out0(inst_cellmath__69), .inst_cellmath__69_0_in0(inst_cellmath__24), .inst_cellmath__69_0_in1(inst_cellmath__19));
cynw_cm_float_cos_inst_cellmath__82_0_bdw1114505291_bdw cynw_cm_float_cos_I19 (.inst_cellmath__82_0_out0(inst_cellmath__82), .inst_cellmath__82_0_in0(inst_cellmath__69), .inst_cellmath__82_0_in1(inst_cellmath__19));
cynw_cm_float_cos_inst_cellmath__66_0_bdw1114505291_bdw cynw_cm_float_cos_I20 (.inst_cellmath__66_0_out0(inst_cellmath__66), .inst_cellmath__66_0_in0(inst_cellmath__24), .inst_cellmath__66_0_in1(inst_cellmath__19), .inst_cellmath__66_0_in2(a_sign));
cynw_cm_float_cos_inst_cellmath__67_0_bdw1114505291_bdw cynw_cm_float_cos_I21 (.inst_cellmath__67_0_out0(inst_cellmath__67), .inst_cellmath__67_0_in0(inst_cellmath__24), .inst_cellmath__67_0_in1(inst_cellmath__19), .inst_cellmath__67_0_in2(a_sign));
cynw_cm_float_cos_inst_cellmath__68_0_bdw1114505291_bdw cynw_cm_float_cos_I22 (.inst_cellmath__68_0_out0(inst_cellmath__68), .inst_cellmath__68_0_in0(inst_cellmath__67), .inst_cellmath__68_0_in1(inst_cellmath__66));
cynw_cm_float_cos_inst_cellmath__228__231__bdw1114505291_bdw cynw_cm_float_cos_I23 (.inst_cellmath__228__231__out0({N741}), .inst_cellmath__228__231__in0({N494}), .inst_cellmath__228__231__in1(inst_cellmath__82), .inst_cellmath__228__231__in2(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__219_0_bdw1114505291_bdw cynw_cm_float_cos_I24 (.inst_cellmath__219_0_out0(inst_cellmath__219), .inst_cellmath__219_0_in0({inst_cellmath__61[22]}), .inst_cellmath__219_0_in1({inst_cellmath__200[48]}));
cynw_cm_float_cos_inst_cellmath__211__182__bdw1114505291_bdw cynw_cm_float_cos_I25 (.inst_cellmath__211__182__out0({N552, N551, N550, N549, N548}), .inst_cellmath__211__182__in0({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_cos_inst_cellmath__215_0_bdw1114505291_bdw cynw_cm_float_cos_I26 (.inst_cellmath__215_0_out0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__215_0_in0({N552, N551, N550, N549, N548}));
cynw_cm_float_cos_inst_cellmath__220__188__bdw1114505291_bdw cynw_cm_float_cos_I27 (.inst_cellmath__220__188__out0({N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661}), .inst_cellmath__220__188__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__220__188__in1({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_cos_inst_cellmath__221__195__bdw1114505291_bdw cynw_cm_float_cos_I28 (.inst_cellmath__221__195__out0({N659, N658, N657, N656, N655, N654, N653}), .inst_cellmath__221__195__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}));
cynw_cm_float_cos_inst_cellmath__220_2WWMM_bdw1114505291_bdw cynw_cm_float_cos_I29 (.inst_cellmath__220_2WWMM_out0({N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709}), .inst_cellmath__220_2WWMM_in0({N659, N658, N657, N656, N655, N654, N653}), .inst_cellmath__220_2WWMM_in1({N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661}), .inst_cellmath__220_2WWMM_in2(inst_cellmath__219));
cynw_cm_float_cos_inst_cellmath__223__208__bdw1114505291_bdw cynw_cm_float_cos_I30 (.inst_cellmath__223__208__out0({N583}), .inst_cellmath__223__208__in0({N715, N714, N713, N712, N711, N710, N709}), .inst_cellmath__223__208__in1({N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717}));
cynw_cm_float_cos_inst_cellmath__223__199__bdw1114505291_bdw cynw_cm_float_cos_I31 (.inst_cellmath__223__199__out0({x[31]}), .inst_cellmath__223__199__in0(inst_cellmath__82), .inst_cellmath__223__199__in1({N493}), .inst_cellmath__223__199__in2({inst_cellmath__42[8], inst_cellmath__42[7], inst_cellmath__42[6]}), .inst_cellmath__223__199__in3({N583}));
cynw_cm_float_cos_inst_cellmath__224__213__bdw1114505291_bdw cynw_cm_float_cos_I32 (.inst_cellmath__224__213__out0({N585}), .inst_cellmath__224__213__in0({N494}), .inst_cellmath__224__213__in1(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__224__212__bdw1114505291_bdw cynw_cm_float_cos_I33 (.inst_cellmath__224__212__out0({N595}), .inst_cellmath__224__212__in0(inst_cellmath__82), .inst_cellmath__224__212__in1({N585}));
cynw_cm_float_cos_inst_cellmath__225__215__bdw1114505291_bdw cynw_cm_float_cos_I34 (.inst_cellmath__225__215__out0({N594}), .inst_cellmath__225__215__in0(inst_cellmath__82), .inst_cellmath__225__215__in1(inst_cellmath__68));
cynw_cm_float_cos_inst_cellmath__228_0_bdw1114505291_bdw cynw_cm_float_cos_I35 (.inst_cellmath__228_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__228_0_in0({N741}), .inst_cellmath__228_0_in1({N594}), .inst_cellmath__228_0_in2({N595}), .inst_cellmath__228_0_in3({N715, N714, N713, N712, N711, N710, N709}));
cynw_cm_float_cos_inst_cellmath__231_0_bdw1114505291_bdw cynw_cm_float_cos_I36 (.inst_cellmath__231_0_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__231_0_in0(inst_cellmath__82), .inst_cellmath__231_0_in1({N741}), .inst_cellmath__231_0_in2({N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717}), .inst_cellmath__231_0_in3({inst_cellmath__210[21]}));
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__200[25] = inst_cellmath__210[0];
assign inst_cellmath__200[26] = inst_cellmath__210[1];
assign inst_cellmath__200[27] = inst_cellmath__210[2];
assign inst_cellmath__200[28] = inst_cellmath__210[3];
assign inst_cellmath__200[29] = inst_cellmath__210[4];
assign inst_cellmath__200[30] = inst_cellmath__210[5];
assign inst_cellmath__200[31] = inst_cellmath__210[6];
assign inst_cellmath__200[32] = inst_cellmath__210[7];
assign inst_cellmath__200[33] = inst_cellmath__210[8];
assign inst_cellmath__200[34] = inst_cellmath__210[9];
assign inst_cellmath__200[35] = inst_cellmath__210[10];
assign inst_cellmath__200[36] = inst_cellmath__210[11];
assign inst_cellmath__200[37] = inst_cellmath__210[12];
assign inst_cellmath__200[38] = inst_cellmath__210[13];
assign inst_cellmath__200[39] = inst_cellmath__210[14];
assign inst_cellmath__200[40] = inst_cellmath__210[15];
assign inst_cellmath__200[41] = inst_cellmath__210[16];
assign inst_cellmath__200[42] = inst_cellmath__210[17];
assign inst_cellmath__200[43] = inst_cellmath__210[18];
assign inst_cellmath__200[44] = inst_cellmath__210[19];
assign inst_cellmath__200[45] = inst_cellmath__210[20];
assign inst_cellmath__200[46] = inst_cellmath__210[21];
assign inst_cellmath__200[47] = inst_cellmath__210[22];
assign inst_cellmath__200[49] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_blk01_cellmath__39_bdw1114505291_bdw (
	inst_blk01_cellmath__39_out0,
	inst_blk01_cellmath__39_in0
	); /* architecture "gate_level" */ 
output [55:0] inst_blk01_cellmath__39_out0;
input [22:0] inst_blk01_cellmath__39_in0;
wire N356,N360,N362,N366,N368,N370,N372 
	,N374,N376,N378,N380,N382,N384,N386,N388 
	,N390,N392,N394,N396,N1066,N1067,N1070,N1071 
	,N1072,N1073,N1078,N1079,N1080,N1081,N1082,N1083 
	,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091 
	,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099 
	,N1100,N1101,N1102,N1103,N1104,N1107,N1108,N1109 
	,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117 
	,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125 
	,N1126,N1127,N1128,N1129,N1132,N1133,N1134,N1135 
	,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143 
	,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151 
	,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159 
	,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167 
	,N1168,N1169,N1170,N1171,N1174,N1175,N1176,N1177 
	,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185 
	,N1186,N1187,N1188,N1189,N1190,N1193,N1194,N1195 
	,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1205 
	,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213 
	,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221 
	,N1222,N1223,N1226,N1227,N1228,N1229,N1230,N1231 
	,N1232,N1233,N1234,N1235,N1238,N1239,N1240,N1241 
	,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249 
	,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257 
	,N1258,N1261,N1262,N1263,N1264,N1265,N1266,N1267 
	,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275 
	,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283 
	,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291 
	,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299 
	,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307 
	,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315 
	,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323 
	,N1324,N1325,N1326,N1327,N1328,N1331,N1332,N1333 
	,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341 
	,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349 
	,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1359 
	,N1360,N1361,N1362,N1363,N1366,N1367,N1368,N1369 
	,N1370,N1373,N1374,N1375,N1376,N1377,N1380,N1381 
	,N1382,N1383,N1384,N1387,N1388,N1389,N1390,N1391 
	,N1392,N1393,N1394,N1395,N1396,N1397,N1404,N1405 
	,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413 
	,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421 
	,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429 
	,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1445 
	,N1446,N1456,N1474,N1476,N1492,N1508,N1528,N1556 
	,N1558,N1562,N1563,N1566,N1567,N1612,N1652,N1654 
	,N1658,N1659,N1694,N1713,N1716,N1719,N1722,N1725 
	,N1728,N1731,N1734,N1737,N1740,N1743,N1746,N1749 
	,N1752,N1755,N1758,N1779,N1782,N1783,N1784,N1786 
	,N1787,N1788,N1790,N1791,N1792,N1794,N1795,N1796 
	,N1798,N1799,N1800,N1802,N1803,N1804,N1806,N1807 
	,N1808,N1810,N1811,N1812,N1814,N1815,N1816,N1818 
	,N1819,N1820,N1822,N1823,N1824,N1826,N1827,N1828 
	,N1830,N1831,N1832,N1834,N1835,N1836,N1838,N1839 
	,N1840,N1842,N1843,N1844,N1846,N1849,N1851,N1852 
	,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860 
	,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868 
	,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876 
	,N1877,N1878,N1879,N1880,N1883,N1885,N1886,N1887 
	,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895 
	,N1896,N1897,N1898,N1899,N1901,N1902,N1905,N1906 
	,N1907,N1910,N1911,N1913,N1914,N1915,N1919,N1923 
	,N1924,N1925,N1927,N1929,N1930,N1931,N1935,N1939 
	,N1940,N1941,N1945,N1949,N1953,N1954,N1955,N1959 
	,N1960,N1961,N1966,N1967,N1969,N1970,N1971,N1975 
	,N1979,N1980,N1981,N1985,N1989,N1993,N1994,N1995 
	,N1999,N2000,N2001,N2005,N2009,N2013,N2017,N2021 
	,N2022,N2023,N2027,N2028,N2029,N2033,N2034,N2035 
	,N2039,N2040,N2041,N2045,N2046,N2047,N2051,N2199 
	,N2212,N2225,N2238,N2251,N2270,N2283,N2296,N2309 
	,N2322,N2341,N2354,N2367,N2380,N2393,N2406,N2419 
	,N2432,N2445,N2458,N2480,N2493,N2506,N2519,N2532 
	,N2554,N2567,N2589,N2602,N2615,N2628,N2641,N2663 
	,N2676,N2698,N2711,N2724,N2737,N2750,N2769,N2782 
	,N2795,N2808,N2821,N2834,N2847,N2860,N2873,N2886 
	,N2899,N2912,N2925,N2938,N2951,N2964,N2983,N2996 
	,N3009,N3022,N3035,N3048,N3067,N3086,N3105,N3124 
	,N3146,N3251,N3254,N3261,N3274,N3282,N3290,N3291 
	,N3305,N3306,N3319,N3333,N3342,N3343,N3361,N3365 
	,N3374,N3375,N3376,N3378,N3379,N3380,N3381,N3382 
	,N3383,N3384,N3385,N3386,N3387,N3388,N3407,N3414 
	,N3441,N3443;
INVXL inst_blk01_cellmath__39_I1377 (.Y(N3251), .A(inst_blk01_cellmath__39_in0[0]));
INVXL inst_blk01_cellmath__39_I1380 (.Y(N3254), .A(inst_blk01_cellmath__39_in0[1]));
INVXL inst_blk01_cellmath__39_I7 (.Y(N356), .A(inst_blk01_cellmath__39_in0[2]));
INVXL inst_blk01_cellmath__39_I8 (.Y(N1067), .A(inst_blk01_cellmath__39_in0[3]));
INVXL inst_blk01_cellmath__39_I9 (.Y(N360), .A(inst_blk01_cellmath__39_in0[4]));
INVXL inst_blk01_cellmath__39_I10 (.Y(N362), .A(inst_blk01_cellmath__39_in0[5]));
INVXL inst_blk01_cellmath__39_I1387 (.Y(N3261), .A(inst_blk01_cellmath__39_in0[6]));
INVXL inst_blk01_cellmath__39_I12 (.Y(N366), .A(inst_blk01_cellmath__39_in0[7]));
INVXL inst_blk01_cellmath__39_I13 (.Y(N368), .A(inst_blk01_cellmath__39_in0[8]));
INVXL inst_blk01_cellmath__39_I14 (.Y(N370), .A(inst_blk01_cellmath__39_in0[9]));
INVXL inst_blk01_cellmath__39_I15 (.Y(N372), .A(inst_blk01_cellmath__39_in0[10]));
INVXL inst_blk01_cellmath__39_I16 (.Y(N374), .A(inst_blk01_cellmath__39_in0[11]));
INVXL inst_blk01_cellmath__39_I17 (.Y(N376), .A(inst_blk01_cellmath__39_in0[12]));
INVXL inst_blk01_cellmath__39_I18 (.Y(N378), .A(inst_blk01_cellmath__39_in0[13]));
INVXL inst_blk01_cellmath__39_I19 (.Y(N380), .A(inst_blk01_cellmath__39_in0[14]));
INVXL inst_blk01_cellmath__39_I20 (.Y(N382), .A(inst_blk01_cellmath__39_in0[15]));
INVXL inst_blk01_cellmath__39_I21 (.Y(N384), .A(inst_blk01_cellmath__39_in0[16]));
INVXL inst_blk01_cellmath__39_I22 (.Y(N386), .A(inst_blk01_cellmath__39_in0[17]));
INVXL inst_blk01_cellmath__39_I23 (.Y(N388), .A(inst_blk01_cellmath__39_in0[18]));
INVXL inst_blk01_cellmath__39_I24 (.Y(N390), .A(inst_blk01_cellmath__39_in0[19]));
INVXL inst_blk01_cellmath__39_I25 (.Y(N392), .A(inst_blk01_cellmath__39_in0[20]));
INVXL inst_blk01_cellmath__39_I26 (.Y(N394), .A(inst_blk01_cellmath__39_in0[21]));
INVXL inst_blk01_cellmath__39_I27 (.Y(N396), .A(inst_blk01_cellmath__39_in0[22]));
INVXL inst_blk01_cellmath__39_I331 (.Y(N1066), .A(N1067));
ADDHX1 inst_blk01_cellmath__39_I332 (.CO(N1071), .S(N1070), .A(N360), .B(N1067));
ADDHX1 inst_blk01_cellmath__39_I333 (.CO(N1073), .S(N1072), .A(N362), .B(N356));
ADDFX1 inst_blk01_cellmath__39_I335 (.CO(N1079), .S(N1078), .A(N3251), .B(N1067), .CI(inst_blk01_cellmath__39_in0[6]));
ADDHX1 inst_blk01_cellmath__39_I336 (.CO(N1081), .S(N1080), .A(N366), .B(N3261));
ADDFX1 inst_blk01_cellmath__39_I337 (.CO(N1083), .S(N1082), .A(N3254), .B(N360), .CI(N1080));
ADDHX1 inst_blk01_cellmath__39_I338 (.CO(N1085), .S(N1084), .A(N368), .B(N362));
ADDFX1 inst_blk01_cellmath__39_I339 (.CO(N1087), .S(N1086), .A(N1081), .B(N356), .CI(N1084));
ADDFX1 arith_dfa_A_I1150 (.CO(N1090), .S(N2199), .A(N3261), .B(inst_blk01_cellmath__39_in0[0]), .CI(N370));
ADDFX1 arith_dfa_A_I1151 (.CO(N1089), .S(N1088), .A(N1067), .B(N1085), .CI(N2199));
ADDFX1 arith_dfa_A_I1152 (.CO(N1093), .S(N2212), .A(N372), .B(inst_blk01_cellmath__39_in0[1]), .CI(N366));
ADDFX1 arith_dfa_A_I1153 (.CO(N1092), .S(N1091), .A(N360), .B(N1090), .CI(N2212));
ADDFX1 arith_dfa_A_I1154 (.CO(N1096), .S(N2225), .A(N368), .B(inst_blk01_cellmath__39_in0[2]), .CI(N374));
ADDFX1 arith_dfa_A_I1155 (.CO(N1095), .S(N1094), .A(N362), .B(N1093), .CI(N2225));
ADDFX1 arith_dfa_A_I1156 (.CO(N1099), .S(N2238), .A(N376), .B(inst_blk01_cellmath__39_in0[3]), .CI(N370));
ADDFX1 arith_dfa_A_I1157 (.CO(N1098), .S(N1097), .A(N1096), .B(N3261), .CI(N2238));
ADDFX1 arith_dfa_A_I1158 (.CO(N1102), .S(N2251), .A(N378), .B(inst_blk01_cellmath__39_in0[4]), .CI(N372));
ADDFX1 arith_dfa_A_I1159 (.CO(N1101), .S(N1100), .A(N366), .B(N1099), .CI(N2251));
XNOR2X1 hap1_A_I1160 (.Y(N1103), .A(inst_blk01_cellmath__39_in0[5]), .B(N3251));
OR2XL hap1_A_I1161 (.Y(N1104), .A(inst_blk01_cellmath__39_in0[5]), .B(N3251));
ADDFX1 arith_dfa_A_I1162 (.CO(N1109), .S(N2270), .A(N374), .B(N380), .CI(N368));
ADDFX1 arith_dfa_A_I1163 (.CO(N1108), .S(N1107), .A(N1102), .B(N1103), .CI(N2270));
ADDFX1 inst_blk01_cellmath__39_I347 (.CO(N1111), .S(N1110), .A(N3254), .B(inst_blk01_cellmath__39_in0[6]), .CI(N382));
ADDFX1 arith_dfa_A_I1164 (.CO(N1114), .S(N2283), .A(N370), .B(N376), .CI(N1104));
ADDFX1 arith_dfa_A_I1165 (.CO(N1113), .S(N1112), .A(N1109), .B(N1110), .CI(N2283));
ADDHX1 inst_blk01_cellmath__39_I349 (.CO(N1116), .S(N1115), .A(inst_blk01_cellmath__39_in0[7]), .B(N356));
ADDFX1 inst_blk01_cellmath__39_I350 (.CO(N1118), .S(N1117), .A(N384), .B(inst_blk01_cellmath__39_in0[0]), .CI(N378));
ADDFX1 arith_dfa_A_I1166 (.CO(N1121), .S(N2296), .A(N1115), .B(N372), .CI(N1111));
ADDFX1 arith_dfa_A_I1167 (.CO(N1120), .S(N1119), .A(N1117), .B(N1114), .CI(N2296));
ADDFX1 arith_dfa_A_I1168 (.CO(N1124), .S(N2309), .A(N1067), .B(inst_blk01_cellmath__39_in0[8]), .CI(N386));
ADDFX1 arith_dfa_A_I1169 (.CO(N1123), .S(N1122), .A(N1116), .B(N1118), .CI(N2309));
ADDFX1 arith_dfa_A_I1170 (.CO(N1127), .S(N2322), .A(N374), .B(inst_blk01_cellmath__39_in0[1]), .CI(N380));
ADDFX1 arith_dfa_A_I1171 (.CO(N1126), .S(N1125), .A(N1122), .B(N1121), .CI(N2322));
XNOR2X1 hap1_A_I1172 (.Y(N1128), .A(inst_blk01_cellmath__39_in0[9]), .B(N360));
OR2XL hap1_A_I1173 (.Y(N1129), .A(inst_blk01_cellmath__39_in0[9]), .B(N360));
ADDFX1 arith_dfa_A_I1174 (.CO(N1134), .S(N2341), .A(N388), .B(inst_blk01_cellmath__39_in0[2]), .CI(N382));
ADDFX1 arith_dfa_A_I1175 (.CO(N1133), .S(N1132), .A(N1127), .B(N1124), .CI(N2341));
ADDFX1 arith_dfa_A_I1176 (.CO(N1137), .S(N2354), .A(N3251), .B(N376), .CI(N1128));
ADDFX1 arith_dfa_A_I1177 (.CO(N1136), .S(N1135), .A(N1132), .B(N1123), .CI(N2354));
ADDFX1 inst_blk01_cellmath__39_I357 (.CO(N1139), .S(N1138), .A(N362), .B(inst_blk01_cellmath__39_in0[10]), .CI(N390));
ADDFX1 arith_dfa_A_I1178 (.CO(N1142), .S(N2367), .A(N384), .B(inst_blk01_cellmath__39_in0[3]), .CI(N378));
ADDFX1 arith_dfa_A_I1179 (.CO(N1141), .S(N1140), .A(N1134), .B(N1138), .CI(N2367));
ADDFX1 arith_dfa_A_I1180 (.CO(N1145), .S(N2380), .A(N1129), .B(N3254), .CI(N1137));
ADDFX1 arith_dfa_A_I1181 (.CO(N1144), .S(N1143), .A(N1133), .B(N1140), .CI(N2380));
ADDFX1 inst_blk01_cellmath__39_I360 (.CO(N1147), .S(N1146), .A(N3261), .B(inst_blk01_cellmath__39_in0[11]), .CI(N392));
ADDFX1 arith_dfa_A_I1182 (.CO(N1150), .S(N2393), .A(N386), .B(inst_blk01_cellmath__39_in0[4]), .CI(N380));
ADDFX1 arith_dfa_A_I1183 (.CO(N1149), .S(N1148), .A(N1142), .B(N1146), .CI(N2393));
ADDFX1 arith_dfa_A_I1184 (.CO(N1153), .S(N2406), .A(N1139), .B(N356), .CI(N1141));
ADDFX1 arith_dfa_A_I1185 (.CO(N1152), .S(N1151), .A(N1145), .B(N1148), .CI(N2406));
ADDFX1 inst_blk01_cellmath__39_I363 (.CO(N1155), .S(N1154), .A(N366), .B(inst_blk01_cellmath__39_in0[12]), .CI(N394));
ADDFX1 arith_dfa_A_I1186 (.CO(N1158), .S(N2419), .A(N382), .B(inst_blk01_cellmath__39_in0[5]), .CI(N388));
ADDFX1 arith_dfa_A_I1187 (.CO(N1157), .S(N1156), .A(N1150), .B(N1154), .CI(N2419));
ADDFX1 arith_dfa_A_I1188 (.CO(N1161), .S(N2432), .A(N1147), .B(N1067), .CI(N1149));
ADDFX1 arith_dfa_A_I1189 (.CO(N1160), .S(N1159), .A(N1156), .B(N1153), .CI(N2432));
ADDFX1 inst_blk01_cellmath__39_I366 (.CO(N1163), .S(N1162), .A(N368), .B(inst_blk01_cellmath__39_in0[13]), .CI(N396));
ADDFX1 arith_dfa_A_I1190 (.CO(N1166), .S(N2445), .A(N390), .B(inst_blk01_cellmath__39_in0[6]), .CI(N384));
ADDFX1 arith_dfa_A_I1191 (.CO(N1165), .S(N1164), .A(N1158), .B(N2445), .CI(N1162));
ADDFX1 arith_dfa_A_I1192 (.CO(N1169), .S(N2458), .A(N1155), .B(N360), .CI(N1157));
ADDFX1 arith_dfa_A_I1193 (.CO(N1168), .S(N1167), .A(N1164), .B(N1161), .CI(N2458));
ADDFX1 inst_blk01_cellmath__39_I1195 (.CO(N1171), .S(N1170), .A(N392), .B(N380), .CI(N370));
ADDFX1 arith_dfa_A_I1196 (.CO(N1176), .S(N2480), .A(N386), .B(inst_blk01_cellmath__39_in0[7]), .CI(N362));
ADDFX1 arith_dfa_A_I1197 (.CO(N1175), .S(N1174), .A(N1163), .B(N1166), .CI(N2480));
ADDFX1 arith_dfa_A_I1198 (.CO(N1179), .S(N2493), .A(N1170), .B(N3251), .CI(N1165));
ADDFX1 arith_dfa_A_I1199 (.CO(N1178), .S(N1177), .A(N1169), .B(N1174), .CI(N2493));
XNOR2X1 hap1_A_I1589 (.Y(N2506), .A(inst_blk01_cellmath__39_in0[15]), .B(N372));
OR2XL hap1_A_I1590 (.Y(N1182), .A(inst_blk01_cellmath__39_in0[15]), .B(N372));
ADDFX1 arith_dfa_A_I1201 (.CO(N1181), .S(N1180), .A(N1176), .B(N1171), .CI(N2506));
ADDFX1 arith_dfa_A_I1202 (.CO(N1185), .S(N2519), .A(N394), .B(inst_blk01_cellmath__39_in0[8]), .CI(N388));
ADDFX1 arith_dfa_A_I1203 (.CO(N1184), .S(N1183), .A(N3254), .B(N3261), .CI(N2519));
ADDFX1 arith_dfa_A_I1204 (.CO(N1188), .S(N2532), .A(N1175), .B(inst_blk01_cellmath__39_in0[14]), .CI(N1180));
ADDFX1 arith_dfa_A_I1205 (.CO(N1187), .S(N1186), .A(N1183), .B(N1179), .CI(N2532));
ADDFX1 inst_blk01_cellmath__39_I1207 (.CO(N1190), .S(N1189), .A(N396), .B(N374), .CI(N384));
ADDFX1 inst_blk01_cellmath__39_I376 (.CO(N1194), .S(N1193), .A(N390), .B(inst_blk01_cellmath__39_in0[9]), .CI(N366));
ADDFX1 arith_dfa_A_I1208 (.CO(N1197), .S(N2554), .A(N356), .B(inst_blk01_cellmath__39_in0[0]), .CI(N1182));
ADDFX1 arith_dfa_A_I1209 (.CO(N1196), .S(N1195), .A(N1193), .B(N1189), .CI(N2554));
ADDFX1 arith_dfa_A_I1210 (.CO(N1200), .S(N2567), .A(N1181), .B(N1185), .CI(N1184));
ADDFX1 arith_dfa_A_I1211 (.CO(N1199), .S(N1198), .A(N1195), .B(N1188), .CI(N2567));
ADDFX1 inst_blk01_cellmath__39_I1213 (.CO(N1202), .S(N1201), .A(N392), .B(N376), .CI(N386));
ADDFX1 inst_blk01_cellmath__39_I380 (.CO(N1206), .S(N1205), .A(N368), .B(inst_blk01_cellmath__39_in0[10]), .CI(N1067));
ADDFX1 arith_dfa_A_I1214 (.CO(N1209), .S(N2589), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[1]), .CI(N1194));
ADDFX1 arith_dfa_A_I1215 (.CO(N1208), .S(N1207), .A(N1201), .B(N1197), .CI(N2589));
ADDFX1 arith_dfa_A_I1216 (.CO(N1212), .S(N2602), .A(N1205), .B(N1190), .CI(N1196));
ADDFX1 arith_dfa_A_I1217 (.CO(N1211), .S(N1210), .A(N1200), .B(N1207), .CI(N2602));
ADDFX1 arith_dfa_A_I1218 (.CO(N1215), .S(N2615), .A(N378), .B(inst_blk01_cellmath__39_in0[18]), .CI(N394));
ADDFX1 arith_dfa_A_I1219 (.CO(N1214), .S(N1213), .A(N1206), .B(N1202), .CI(N2615));
ADDFX1 arith_dfa_A_I1220 (.CO(N1218), .S(N2628), .A(N360), .B(inst_blk01_cellmath__39_in0[11]), .CI(N370));
ADDFX1 arith_dfa_A_I1221 (.CO(N1217), .S(N1216), .A(inst_blk01_cellmath__39_in0[17]), .B(inst_blk01_cellmath__39_in0[2]), .CI(N2628));
ADDFX1 arith_dfa_A_I1222 (.CO(N1221), .S(N2641), .A(N1213), .B(N1209), .CI(N1216));
ADDFX1 arith_dfa_A_I1223 (.CO(N1220), .S(N1219), .A(N1208), .B(N1212), .CI(N2641));
ADDFX1 inst_blk01_cellmath__39_I1225 (.CO(N1223), .S(N1222), .A(N396), .B(N380), .CI(N390));
ADDFX1 inst_blk01_cellmath__39_I387 (.CO(N1227), .S(N1226), .A(N372), .B(inst_blk01_cellmath__39_in0[12]), .CI(N362));
ADDFX1 arith_dfa_A_I1226 (.CO(N1230), .S(N2663), .A(inst_blk01_cellmath__39_in0[0]), .B(inst_blk01_cellmath__39_in0[3]), .CI(N1215));
ADDFX1 arith_dfa_A_I1227 (.CO(N1229), .S(N1228), .A(N1226), .B(N1222), .CI(N2663));
ADDFX1 arith_dfa_A_I1228 (.CO(N1233), .S(N2676), .A(N1214), .B(N1218), .CI(N1217));
ADDFX1 arith_dfa_A_I1229 (.CO(N1232), .S(N1231), .A(N1221), .B(N1228), .CI(N2676));
ADDFX1 inst_blk01_cellmath__39_I1231 (.CO(N1235), .S(N1234), .A(N374), .B(N382), .CI(N392));
ADDFX1 inst_blk01_cellmath__39_I391 (.CO(N1239), .S(N1238), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[13]), .CI(N3261));
ADDFX1 arith_dfa_A_I1232 (.CO(N1242), .S(N2698), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[1]), .CI(N1227));
ADDFX1 arith_dfa_A_I1233 (.CO(N1241), .S(N1240), .A(N1234), .B(N1230), .CI(N2698));
ADDFX1 arith_dfa_A_I1234 (.CO(N1245), .S(N2711), .A(N1238), .B(N1223), .CI(N1229));
ADDFX1 arith_dfa_A_I1235 (.CO(N1244), .S(N1243), .A(N1233), .B(N1240), .CI(N2711));
ADDHX1 inst_blk01_cellmath__39_I394 (.CO(N1247), .S(N1246), .A(inst_blk01_cellmath__39_in0[21]), .B(N384));
ADDFX1 arith_dfa_A_I1236 (.CO(N1250), .S(N2724), .A(N376), .B(inst_blk01_cellmath__39_in0[14]), .CI(N366));
ADDFX1 arith_dfa_A_I1237 (.CO(N1249), .S(N1248), .A(N1239), .B(N1235), .CI(N2724));
ADDFX1 arith_dfa_A_I1238 (.CO(N1253), .S(N2737), .A(inst_blk01_cellmath__39_in0[2]), .B(inst_blk01_cellmath__39_in0[5]), .CI(inst_blk01_cellmath__39_in0[0]));
ADDFX1 arith_dfa_A_I1239 (.CO(N1252), .S(N1251), .A(inst_blk01_cellmath__39_in0[20]), .B(N1246), .CI(N2737));
ADDFX1 arith_dfa_A_I1240 (.CO(N1256), .S(N2750), .A(N1251), .B(N1242), .CI(N1248));
ADDFX1 arith_dfa_A_I1241 (.CO(N1255), .S(N1254), .A(N1241), .B(N1245), .CI(N2750));
XNOR2X1 hap1_A_I1242 (.Y(N1257), .A(N386), .B(N378));
OR2XL hap1_A_I1243 (.Y(N1258), .A(N386), .B(N378));
ADDFX1 arith_dfa_A_I1244 (.CO(N1263), .S(N2769), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[22]), .CI(N368));
ADDFX1 arith_dfa_A_I1245 (.CO(N1262), .S(N1261), .A(N1250), .B(N1257), .CI(N2769));
ADDFX1 arith_dfa_A_I1246 (.CO(N1266), .S(N2782), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[6]), .CI(inst_blk01_cellmath__39_in0[1]));
ADDFX1 arith_dfa_A_I1247 (.CO(N1265), .S(N1264), .A(N1247), .B(N1253), .CI(N2782));
ADDFX1 arith_dfa_A_I1248 (.CO(N1269), .S(N2795), .A(N1249), .B(N1252), .CI(N1264));
ADDFX1 arith_dfa_A_I1249 (.CO(N1268), .S(N1267), .A(N1261), .B(N1256), .CI(N2795));
ADDFX1 arith_dfa_A_I1250 (.CO(N1272), .S(N2808), .A(N388), .B(inst_blk01_cellmath__39_in0[16]), .CI(N380));
ADDFX1 arith_dfa_A_I1251 (.CO(N1271), .S(N1270), .A(N1266), .B(N1263), .CI(N2808));
ADDFX1 arith_dfa_A_I1252 (.CO(N1275), .S(N2821), .A(N370), .B(inst_blk01_cellmath__39_in0[7]), .CI(inst_blk01_cellmath__39_in0[4]));
ADDFX1 arith_dfa_A_I1253 (.CO(N1274), .S(N1273), .A(inst_blk01_cellmath__39_in0[2]), .B(N1258), .CI(N2821));
ADDFX1 arith_dfa_A_I1254 (.CO(N1278), .S(N2834), .A(N1262), .B(N1265), .CI(N1270));
ADDFX1 arith_dfa_A_I1255 (.CO(N1277), .S(N1276), .A(N1273), .B(N1269), .CI(N2834));
ADDHX1 inst_blk01_cellmath__39_I405 (.CO(N1280), .S(N1279), .A(inst_blk01_cellmath__39_in0[17]), .B(N390));
ADDFX1 inst_blk01_cellmath__39_I406 (.CO(N1282), .S(N1281), .A(N382), .B(inst_blk01_cellmath__39_in0[8]), .CI(N372));
ADDFX1 arith_dfa_A_I1256 (.CO(N1285), .S(N2847), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[5]), .CI(N1279));
ADDFX1 arith_dfa_A_I1257 (.CO(N1284), .S(N1283), .A(N1272), .B(N1281), .CI(N2847));
ADDFX1 arith_dfa_A_I1258 (.CO(N1288), .S(N2860), .A(N1271), .B(N1275), .CI(N1274));
ADDFX1 arith_dfa_A_I1259 (.CO(N1287), .S(N1286), .A(N1278), .B(N1283), .CI(N2860));
ADDHX1 inst_blk01_cellmath__39_I409 (.CO(N1290), .S(N1289), .A(inst_blk01_cellmath__39_in0[18]), .B(N392));
ADDFX1 inst_blk01_cellmath__39_I410 (.CO(N1292), .S(N1291), .A(N384), .B(inst_blk01_cellmath__39_in0[9]), .CI(N374));
ADDFX1 arith_dfa_A_I1260 (.CO(N1295), .S(N2873), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[6]), .CI(N1280));
ADDFX1 arith_dfa_A_I1261 (.CO(N1294), .S(N1293), .A(N1291), .B(N1285), .CI(N2873));
ADDFX1 arith_dfa_A_I1262 (.CO(N1298), .S(N2886), .A(N1282), .B(N1289), .CI(N1284));
ADDFX1 arith_dfa_A_I1263 (.CO(N1297), .S(N1296), .A(N1293), .B(N1288), .CI(N2886));
ADDHX1 inst_blk01_cellmath__39_I413 (.CO(N1300), .S(N1299), .A(inst_blk01_cellmath__39_in0[19]), .B(N394));
ADDFX1 inst_blk01_cellmath__39_I414 (.CO(N1302), .S(N1301), .A(N386), .B(inst_blk01_cellmath__39_in0[10]), .CI(N376));
ADDFX1 arith_dfa_A_I1264 (.CO(N1305), .S(N2899), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[7]), .CI(N1290));
ADDFX1 arith_dfa_A_I1265 (.CO(N1304), .S(N1303), .A(N1301), .B(N1295), .CI(N2899));
ADDFX1 arith_dfa_A_I1266 (.CO(N1308), .S(N2912), .A(N1292), .B(N1299), .CI(N1294));
ADDFX1 arith_dfa_A_I1267 (.CO(N1307), .S(N1306), .A(N1303), .B(N1298), .CI(N2912));
ADDHX1 inst_blk01_cellmath__39_I417 (.CO(N1310), .S(N1309), .A(inst_blk01_cellmath__39_in0[20]), .B(N396));
ADDFX1 inst_blk01_cellmath__39_I418 (.CO(N1312), .S(N1311), .A(N388), .B(inst_blk01_cellmath__39_in0[11]), .CI(N378));
ADDFX1 arith_dfa_A_I1268 (.CO(N1315), .S(N2925), .A(inst_blk01_cellmath__39_in0[6]), .B(inst_blk01_cellmath__39_in0[8]), .CI(N1300));
ADDFX1 arith_dfa_A_I1269 (.CO(N1314), .S(N1313), .A(N1311), .B(N1305), .CI(N2925));
ADDFX1 arith_dfa_A_I1270 (.CO(N1318), .S(N2938), .A(N1302), .B(N1309), .CI(N1304));
ADDFX1 arith_dfa_A_I1271 (.CO(N1317), .S(N1316), .A(N1313), .B(N1308), .CI(N2938));
ADDFX1 inst_blk01_cellmath__39_I421 (.CO(N1320), .S(N1319), .A(N390), .B(inst_blk01_cellmath__39_in0[21]), .CI(N380));
ADDFX1 arith_dfa_A_I1272 (.CO(N1323), .S(N2951), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[12]), .CI(inst_blk01_cellmath__39_in0[7]));
ADDFX1 arith_dfa_A_I1273 (.CO(N1322), .S(N1321), .A(N1319), .B(N1315), .CI(N2951));
ADDFX1 arith_dfa_A_I1274 (.CO(N1326), .S(N2964), .A(N1312), .B(N1310), .CI(N1314));
ADDFX1 arith_dfa_A_I1275 (.CO(N1325), .S(N1324), .A(N1321), .B(N1318), .CI(N2964));
XNOR2X1 hap1_A_I1276 (.Y(N1327), .A(N392), .B(N382));
OR2XL hap1_A_I1277 (.Y(N1328), .A(N392), .B(N382));
ADDFX1 arith_dfa_A_I1278 (.CO(N1333), .S(N2983), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[22]), .CI(inst_blk01_cellmath__39_in0[10]));
ADDFX1 arith_dfa_A_I1279 (.CO(N1332), .S(N1331), .A(N1320), .B(N1327), .CI(N2983));
ADDFX1 arith_dfa_A_I1280 (.CO(N1336), .S(N2996), .A(N1323), .B(inst_blk01_cellmath__39_in0[8]), .CI(N1322));
ADDFX1 arith_dfa_A_I1281 (.CO(N1335), .S(N1334), .A(N1331), .B(N1326), .CI(N2996));
ADDFX1 arith_dfa_A_I1282 (.CO(N1339), .S(N3009), .A(N394), .B(inst_blk01_cellmath__39_in0[14]), .CI(N384));
ADDFX1 arith_dfa_A_I1283 (.CO(N1338), .S(N1337), .A(N1328), .B(N1333), .CI(N3009));
ADDFX1 arith_dfa_A_I1284 (.CO(N1342), .S(N3022), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[11]), .CI(N1332));
ADDFX1 arith_dfa_A_I1285 (.CO(N1341), .S(N1340), .A(N1337), .B(N1336), .CI(N3022));
ADDHX1 inst_blk01_cellmath__39_I429 (.CO(N1344), .S(N1343), .A(inst_blk01_cellmath__39_in0[15]), .B(N396));
ADDFX1 inst_blk01_cellmath__39_I430 (.CO(N1346), .S(N1345), .A(inst_blk01_cellmath__39_in0[10]), .B(inst_blk01_cellmath__39_in0[12]), .CI(N386));
ADDFX1 arith_dfa_A_I1286 (.CO(N1349), .S(N3035), .A(N1339), .B(N1343), .CI(N1345));
ADDFX1 arith_dfa_A_I1287 (.CO(N1348), .S(N1347), .A(N1342), .B(N1338), .CI(N3035));
ADDFX1 inst_blk01_cellmath__39_I432 (.CO(N1351), .S(N1350), .A(N388), .B(inst_blk01_cellmath__39_in0[16]), .CI(inst_blk01_cellmath__39_in0[13]));
ADDFX1 arith_dfa_A_I1288 (.CO(N1354), .S(N3048), .A(N1346), .B(inst_blk01_cellmath__39_in0[11]), .CI(N1344));
ADDFX1 arith_dfa_A_I1289 (.CO(N1353), .S(N1352), .A(N1350), .B(N1349), .CI(N3048));
XNOR2X1 hap1_A_I1290 (.Y(N1355), .A(N390), .B(inst_blk01_cellmath__39_in0[17]));
OR2XL hap1_A_I1291 (.Y(N1356), .A(N390), .B(inst_blk01_cellmath__39_in0[17]));
ADDFX1 arith_dfa_A_I1292 (.CO(N1361), .S(N3067), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[14]), .CI(N1351));
ADDFX1 arith_dfa_A_I1293 (.CO(N1360), .S(N1359), .A(N1355), .B(N1354), .CI(N3067));
XNOR2X1 hap1_A_I1294 (.Y(N1362), .A(N392), .B(inst_blk01_cellmath__39_in0[18]));
OR2XL hap1_A_I1295 (.Y(N1363), .A(N392), .B(inst_blk01_cellmath__39_in0[18]));
ADDFX1 arith_dfa_A_I1296 (.CO(N1368), .S(N3086), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[15]), .CI(N1356));
ADDFX1 arith_dfa_A_I1297 (.CO(N1367), .S(N1366), .A(N1362), .B(N1361), .CI(N3086));
XNOR2X1 hap1_A_I1298 (.Y(N1369), .A(N394), .B(inst_blk01_cellmath__39_in0[19]));
OR2XL hap1_A_I1299 (.Y(N1370), .A(N394), .B(inst_blk01_cellmath__39_in0[19]));
ADDFX1 arith_dfa_A_I1300 (.CO(N1375), .S(N3105), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[16]), .CI(N1363));
ADDFX1 arith_dfa_A_I1301 (.CO(N1374), .S(N1373), .A(N1369), .B(N1368), .CI(N3105));
XNOR2X1 hap1_A_I1302 (.Y(N1376), .A(N396), .B(inst_blk01_cellmath__39_in0[20]));
OR2XL hap1_A_I1303 (.Y(N1377), .A(N396), .B(inst_blk01_cellmath__39_in0[20]));
ADDFX1 arith_dfa_A_I1304 (.CO(N1382), .S(N3124), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[17]), .CI(N1370));
ADDFX1 arith_dfa_A_I1305 (.CO(N1381), .S(N1380), .A(N1376), .B(N1375), .CI(N3124));
ADDFX1 inst_blk01_cellmath__39_I1307 (.CO(N1384), .S(N1383), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[18]), .CI(N394));
ADDFX1 inst_blk01_cellmath__39_I443 (.CO(N1388), .S(N1387), .A(N1382), .B(N1377), .CI(N1383));
ADDFX1 arith_dfa_A_I1308 (.CO(N1391), .S(N3146), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[22]), .CI(inst_blk01_cellmath__39_in0[17]));
ADDFX1 arith_dfa_A_I1309 (.CO(N1390), .S(N1389), .A(inst_blk01_cellmath__39_in0[21]), .B(N1384), .CI(N3146));
ADDFX1 inst_blk01_cellmath__39_I445 (.CO(N1393), .S(N1392), .A(inst_blk01_cellmath__39_in0[18]), .B(inst_blk01_cellmath__39_in0[20]), .CI(N1391));
ADDHX1 inst_blk01_cellmath__39_I446 (.CO(N1395), .S(N1394), .A(inst_blk01_cellmath__39_in0[21]), .B(inst_blk01_cellmath__39_in0[19]));
ADDHX1 inst_blk01_cellmath__39_I447 (.CO(N1397), .S(N1396), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[20]));
INVXL inst_blk01_cellmath__39_I451 (.Y(N1404), .A(N356));
NOR2XL inst_blk01_cellmath__39_I452 (.Y(N1405), .A(N3251), .B(N1066));
NAND2XL inst_blk01_cellmath__39_I453 (.Y(N1406), .A(N3251), .B(N1066));
NOR2XL inst_blk01_cellmath__39_I454 (.Y(N1407), .A(N3254), .B(N1070));
NAND2XL inst_blk01_cellmath__39_I455 (.Y(N1408), .A(N3254), .B(N1070));
NOR2XL inst_blk01_cellmath__39_I1564 (.Y(N1409), .A(N1072), .B(N1071));
NAND2XL inst_blk01_cellmath__39_I457 (.Y(N1410), .A(N1071), .B(N1072));
NOR2XL inst_blk01_cellmath__39_I458 (.Y(N1411), .A(N1073), .B(N1078));
NAND2XL inst_blk01_cellmath__39_I459 (.Y(N1412), .A(N1073), .B(N1078));
NOR2XL inst_blk01_cellmath__39_I460 (.Y(N1413), .A(N1079), .B(N1082));
NAND2XL inst_blk01_cellmath__39_I461 (.Y(N1414), .A(N1079), .B(N1082));
NOR2XL inst_blk01_cellmath__39_I462 (.Y(N1415), .A(N1083), .B(N1086));
NAND2XL inst_blk01_cellmath__39_I463 (.Y(N1416), .A(N1083), .B(N1086));
NOR2XL inst_blk01_cellmath__39_I464 (.Y(N1417), .A(N1087), .B(N1088));
NAND2XL inst_blk01_cellmath__39_I465 (.Y(N1418), .A(N1087), .B(N1088));
NOR2XL inst_blk01_cellmath__39_I466 (.Y(N1419), .A(N1089), .B(N1091));
NAND2XL inst_blk01_cellmath__39_I467 (.Y(N1420), .A(N1089), .B(N1091));
NOR2XL inst_blk01_cellmath__39_I468 (.Y(N1421), .A(N1092), .B(N1094));
NAND2XL inst_blk01_cellmath__39_I469 (.Y(N1422), .A(N1092), .B(N1094));
NOR2XL inst_blk01_cellmath__39_I470 (.Y(N1423), .A(N1095), .B(N1097));
NAND2XL inst_blk01_cellmath__39_I471 (.Y(N1424), .A(N1095), .B(N1097));
NOR2XL inst_blk01_cellmath__39_I472 (.Y(N1425), .A(N1098), .B(N1100));
NAND2XL inst_blk01_cellmath__39_I473 (.Y(N1426), .A(N1098), .B(N1100));
NOR2XL inst_blk01_cellmath__39_I474 (.Y(N1427), .A(N1101), .B(N1107));
NAND2XL inst_blk01_cellmath__39_I475 (.Y(N1428), .A(N1101), .B(N1107));
NOR2XL inst_blk01_cellmath__39_I476 (.Y(N1429), .A(N1108), .B(N1112));
NAND2XL inst_blk01_cellmath__39_I477 (.Y(N1430), .A(N1108), .B(N1112));
NOR2XL inst_blk01_cellmath__39_I478 (.Y(N1431), .A(N1113), .B(N1119));
NAND2XL inst_blk01_cellmath__39_I479 (.Y(N1432), .A(N1113), .B(N1119));
NOR2XL inst_blk01_cellmath__39_I480 (.Y(N1433), .A(N1120), .B(N1125));
NAND2XL inst_blk01_cellmath__39_I481 (.Y(N1434), .A(N1120), .B(N1125));
NOR2XL inst_blk01_cellmath__39_I482 (.Y(N1435), .A(N1126), .B(N1135));
NAND2XL inst_blk01_cellmath__39_I483 (.Y(N1436), .A(N1126), .B(N1135));
NOR2XL inst_blk01_cellmath__39_I1530 (.Y(N3274), .A(inst_blk01_cellmath__39_in0[1]), .B(inst_blk01_cellmath__39_in0[0]));
AOI21XL inst_blk01_cellmath__39_I490 (.Y(N1445), .A0(N1406), .A1(N1404), .B0(N1405));
INVXL inst_blk01_cellmath__39_I491 (.Y(N1446), .A(N1406));
OAI21XL inst_blk01_cellmath__39_I498 (.Y(N1456), .A0(N1446), .A1(N3274), .B0(N1445));
AO21XL inst_blk01_cellmath__39_I1582 (.Y(N3282), .A0(N1410), .A1(N1407), .B0(N1409));
AOI21XL inst_blk01_cellmath__39_I516 (.Y(N1474), .A0(N1408), .A1(N1456), .B0(N1407));
AOI31X1 inst_blk01_cellmath__39_I2686 (.Y(N1476), .A0(N1410), .A1(N1408), .A2(N1456), .B0(N3282));
INVXL inst_blk01_cellmath__39_I1416 (.Y(N3290), .A(N1411));
INVXL inst_blk01_cellmath__39_I1417 (.Y(N3291), .A(N1412));
OAI21XL inst_blk01_cellmath__39_I534 (.Y(N1492), .A0(N3291), .A1(N1476), .B0(N3290));
AOI21XL inst_blk01_cellmath__39_I550 (.Y(N1508), .A0(N1414), .A1(N1492), .B0(N1413));
INVXL inst_blk01_cellmath__39_I1431 (.Y(N3305), .A(N1415));
INVXL inst_blk01_cellmath__39_I1432 (.Y(N3306), .A(N1416));
OAI21XL inst_blk01_cellmath__39_I570 (.Y(N1528), .A0(N3306), .A1(N1508), .B0(N3305));
AO21XL inst_blk01_cellmath__39_I1535 (.Y(N3319), .A0(N1420), .A1(N1417), .B0(N1419));
AOI21XL inst_blk01_cellmath__39_I598 (.Y(N1556), .A0(N1418), .A1(N1528), .B0(N1417));
AOI31X1 inst_blk01_cellmath__39_I2687 (.Y(N1558), .A0(N1420), .A1(N1418), .A2(N1528), .B0(N3319));
AOI21XL inst_blk01_cellmath__39_I604 (.Y(N1562), .A0(N1424), .A1(N1421), .B0(N1423));
NAND2XL inst_blk01_cellmath__39_I605 (.Y(N1563), .A(N1424), .B(N1422));
INVXL inst_blk01_cellmath__39_I1459 (.Y(N3333), .A(N1426));
AOI21XL inst_blk01_cellmath__39_I608 (.Y(N1566), .A0(N1428), .A1(N1425), .B0(N1427));
NAND2XL inst_blk01_cellmath__39_I609 (.Y(N1567), .A(N1428), .B(N1426));
NOR2XL andori2bb1_A_I1591 (.Y(N3407), .A(N3333), .B(N1562));
NOR2XL andori2bb1_A_I1592 (.Y(N3342), .A(N3407), .B(N1425));
OR2XL inst_blk01_cellmath__39_I1539 (.Y(N3343), .A(N3333), .B(N1563));
OAI21XL orandi31_A_I2688 (.Y(N3443), .A0(N1567), .A1(N1562), .B0(N1566));
NOR3XL orandi31_A_I1602 (.Y(N3441), .A(N1567), .B(N1563), .C(N1558));
OR2XL orandi31_A_I1603 (.Y(N1612), .A(N3441), .B(N3443));
AO21XL inst_blk01_cellmath__39_I1544 (.Y(N3361), .A0(N1432), .A1(N1429), .B0(N1431));
NOR2BX1 inst_blk01_cellmath__39_I1546 (.Y(N3365), .AN(N3274), .B(N1404));
NOR2BX1 andori2bb1_A_I2689 (.Y(N3414), .AN(N1422), .B(N1558));
NOR2XL andori2bb1_A_I1594 (.Y(N3374), .A(N3414), .B(N1421));
OA21X1 inst_blk01_cellmath__39_I1548 (.Y(N3375), .A0(N1563), .A1(N1558), .B0(N1562));
OA21X1 inst_blk01_cellmath__39_I1549 (.Y(N3376), .A0(N3343), .A1(N1558), .B0(N3342));
AOI21XL inst_blk01_cellmath__39_I694 (.Y(N1652), .A0(N1430), .A1(N1612), .B0(N1429));
AOI31X1 inst_blk01_cellmath__39_I2690 (.Y(N1654), .A0(N1432), .A1(N1430), .A2(N1612), .B0(N3361));
INVXL inst_blk01_cellmath__39_I1504 (.Y(N3378), .A(N1433));
INVXL inst_blk01_cellmath__39_I1505 (.Y(N3379), .A(N1434));
AOI21XL inst_blk01_cellmath__39_I700 (.Y(N1658), .A0(N1436), .A1(N1433), .B0(N1435));
NAND2XL inst_blk01_cellmath__39_I701 (.Y(N1659), .A(N1436), .B(N1434));
OAI21XL inst_blk01_cellmath__39_I736 (.Y(N1694), .A0(N3379), .A1(N1654), .B0(N3378));
OAI21XL inst_blk01_cellmath__39_I738 (.Y(N1779), .A0(N1659), .A1(N1654), .B0(N1658));
NAND2BXL inst_blk01_cellmath__39_I751 (.Y(N1713), .AN(N1405), .B(N1406));
NAND2BXL inst_blk01_cellmath__39_I754 (.Y(N1716), .AN(N1407), .B(N1408));
NAND2BXL inst_blk01_cellmath__39_I757 (.Y(N1719), .AN(N1409), .B(N1410));
NAND2BXL inst_blk01_cellmath__39_I760 (.Y(N1722), .AN(N1411), .B(N1412));
NAND2BXL inst_blk01_cellmath__39_I763 (.Y(N1725), .AN(N1413), .B(N1414));
NAND2BXL inst_blk01_cellmath__39_I766 (.Y(N1728), .AN(N1415), .B(N1416));
NAND2BXL inst_blk01_cellmath__39_I769 (.Y(N1731), .AN(N1417), .B(N1418));
NAND2BXL inst_blk01_cellmath__39_I772 (.Y(N1734), .AN(N1419), .B(N1420));
NAND2BXL inst_blk01_cellmath__39_I775 (.Y(N1737), .AN(N1421), .B(N1422));
NAND2BXL inst_blk01_cellmath__39_I778 (.Y(N1740), .AN(N1423), .B(N1424));
NAND2BXL inst_blk01_cellmath__39_I781 (.Y(N1743), .AN(N1425), .B(N1426));
NAND2BXL inst_blk01_cellmath__39_I784 (.Y(N1746), .AN(N1427), .B(N1428));
NAND2BXL inst_blk01_cellmath__39_I787 (.Y(N1749), .AN(N1429), .B(N1430));
NAND2BXL inst_blk01_cellmath__39_I790 (.Y(N1752), .AN(N1431), .B(N1432));
NAND2BXL inst_blk01_cellmath__39_I793 (.Y(N1755), .AN(N1433), .B(N1434));
NAND2BXL inst_blk01_cellmath__39_I796 (.Y(N1758), .AN(N1435), .B(N1436));
XNOR2X1 inst_blk01_cellmath__39_I1339 (.Y(inst_blk01_cellmath__39_out0[2]), .A(N3251), .B(inst_blk01_cellmath__39_in0[1]));
XNOR2X1 inst_blk01_cellmath__39_I1551 (.Y(inst_blk01_cellmath__39_out0[3]), .A(N3274), .B(N1404));
XNOR2X1 inst_blk01_cellmath__39_I800 (.Y(inst_blk01_cellmath__39_out0[4]), .A(N3365), .B(N1713));
XOR2XL inst_blk01_cellmath__39_I1572 (.Y(inst_blk01_cellmath__39_out0[5]), .A(N1456), .B(N1716));
XNOR2X1 inst_blk01_cellmath__39_I1342 (.Y(inst_blk01_cellmath__39_out0[6]), .A(N1474), .B(N1719));
XNOR2X1 inst_blk01_cellmath__39_I1343 (.Y(inst_blk01_cellmath__39_out0[7]), .A(N1476), .B(N1722));
XOR2XL inst_blk01_cellmath__39_I1553 (.Y(inst_blk01_cellmath__39_out0[8]), .A(N1492), .B(N1725));
XNOR2X1 inst_blk01_cellmath__39_I1345 (.Y(inst_blk01_cellmath__39_out0[9]), .A(N1508), .B(N1728));
XOR2XL inst_blk01_cellmath__39_I1554 (.Y(inst_blk01_cellmath__39_out0[10]), .A(N1528), .B(N1731));
XNOR2X1 inst_blk01_cellmath__39_I1347 (.Y(inst_blk01_cellmath__39_out0[11]), .A(N1556), .B(N1734));
XNOR2X1 inst_blk01_cellmath__39_I1348 (.Y(inst_blk01_cellmath__39_out0[12]), .A(N1558), .B(N1737));
XNOR2X1 inst_blk01_cellmath__39_I2691 (.Y(inst_blk01_cellmath__39_out0[13]), .A(N3374), .B(N1740));
XNOR2X1 inst_blk01_cellmath__39_I2692 (.Y(inst_blk01_cellmath__39_out0[14]), .A(N3375), .B(N1743));
XNOR2X1 inst_blk01_cellmath__39_I2693 (.Y(inst_blk01_cellmath__39_out0[15]), .A(N3376), .B(N1746));
XOR2XL inst_blk01_cellmath__39_I1555 (.Y(inst_blk01_cellmath__39_out0[16]), .A(N1612), .B(N1749));
XNOR2X1 inst_blk01_cellmath__39_I813 (.Y(inst_blk01_cellmath__39_out0[17]), .A(N1652), .B(N1752));
XNOR2X1 inst_blk01_cellmath__39_I814 (.Y(inst_blk01_cellmath__39_out0[18]), .A(N1654), .B(N1755));
XOR2XL inst_blk01_cellmath__39_I815 (.Y(inst_blk01_cellmath__39_out0[19]), .A(N1694), .B(N1758));
XOR2XL inst_blk01_cellmath__39_I819 (.Y(N1782), .A(N1136), .B(N1143));
NOR2XL inst_blk01_cellmath__39_I820 (.Y(N1783), .A(N1144), .B(N1151));
XOR2XL inst_blk01_cellmath__39_I821 (.Y(N1784), .A(N1144), .B(N1151));
XOR2XL inst_blk01_cellmath__39_I823 (.Y(N1786), .A(N1152), .B(N1159));
NOR2XL inst_blk01_cellmath__39_I824 (.Y(N1787), .A(N1160), .B(N1167));
XOR2XL inst_blk01_cellmath__39_I825 (.Y(N1788), .A(N1160), .B(N1167));
XOR2XL inst_blk01_cellmath__39_I827 (.Y(N1790), .A(N1168), .B(N1177));
NOR2XL inst_blk01_cellmath__39_I828 (.Y(N1791), .A(N1178), .B(N1186));
XOR2XL inst_blk01_cellmath__39_I829 (.Y(N1792), .A(N1178), .B(N1186));
XOR2XL inst_blk01_cellmath__39_I831 (.Y(N1794), .A(N1187), .B(N1198));
NOR2XL inst_blk01_cellmath__39_I832 (.Y(N1795), .A(N1199), .B(N1210));
XOR2XL inst_blk01_cellmath__39_I833 (.Y(N1796), .A(N1199), .B(N1210));
XOR2XL inst_blk01_cellmath__39_I835 (.Y(N1798), .A(N1211), .B(N1219));
NOR2XL inst_blk01_cellmath__39_I836 (.Y(N1799), .A(N1220), .B(N1231));
XOR2XL inst_blk01_cellmath__39_I837 (.Y(N1800), .A(N1220), .B(N1231));
XOR2XL inst_blk01_cellmath__39_I839 (.Y(N1802), .A(N1232), .B(N1243));
NOR2XL inst_blk01_cellmath__39_I840 (.Y(N1803), .A(N1244), .B(N1254));
XOR2XL inst_blk01_cellmath__39_I841 (.Y(N1804), .A(N1244), .B(N1254));
XOR2XL inst_blk01_cellmath__39_I843 (.Y(N1806), .A(N1255), .B(N1267));
NOR2XL inst_blk01_cellmath__39_I844 (.Y(N1807), .A(N1268), .B(N1276));
XOR2XL inst_blk01_cellmath__39_I845 (.Y(N1808), .A(N1268), .B(N1276));
XOR2XL inst_blk01_cellmath__39_I847 (.Y(N1810), .A(N1277), .B(N1286));
NOR2XL inst_blk01_cellmath__39_I848 (.Y(N1811), .A(N1287), .B(N1296));
XOR2XL inst_blk01_cellmath__39_I849 (.Y(N1812), .A(N1287), .B(N1296));
XOR2XL inst_blk01_cellmath__39_I851 (.Y(N1814), .A(N1297), .B(N1306));
NOR2XL inst_blk01_cellmath__39_I852 (.Y(N1815), .A(N1307), .B(N1316));
XOR2XL inst_blk01_cellmath__39_I853 (.Y(N1816), .A(N1307), .B(N1316));
XOR2XL inst_blk01_cellmath__39_I855 (.Y(N1818), .A(N1317), .B(N1324));
NOR2XL inst_blk01_cellmath__39_I856 (.Y(N1819), .A(N1325), .B(N1334));
XOR2XL inst_blk01_cellmath__39_I857 (.Y(N1820), .A(N1325), .B(N1334));
XOR2XL inst_blk01_cellmath__39_I859 (.Y(N1822), .A(N1335), .B(N1340));
NOR2XL inst_blk01_cellmath__39_I860 (.Y(N1823), .A(N1341), .B(N1347));
XOR2XL inst_blk01_cellmath__39_I861 (.Y(N1824), .A(N1341), .B(N1347));
XOR2XL inst_blk01_cellmath__39_I863 (.Y(N1826), .A(N1352), .B(N1348));
NOR2XL inst_blk01_cellmath__39_I864 (.Y(N1827), .A(N1353), .B(N1359));
XOR2XL inst_blk01_cellmath__39_I865 (.Y(N1828), .A(N1353), .B(N1359));
XOR2XL inst_blk01_cellmath__39_I867 (.Y(N1830), .A(N1360), .B(N1366));
NOR2XL inst_blk01_cellmath__39_I868 (.Y(N1831), .A(N1367), .B(N1373));
XOR2XL inst_blk01_cellmath__39_I869 (.Y(N1832), .A(N1367), .B(N1373));
XOR2XL inst_blk01_cellmath__39_I871 (.Y(N1834), .A(N1374), .B(N1380));
NOR2XL inst_blk01_cellmath__39_I872 (.Y(N1835), .A(N1387), .B(N1381));
XOR2XL inst_blk01_cellmath__39_I873 (.Y(N1836), .A(N1387), .B(N1381));
XOR2XL inst_blk01_cellmath__39_I875 (.Y(N1838), .A(N1388), .B(N1389));
NOR2XL inst_blk01_cellmath__39_I876 (.Y(N1839), .A(N1392), .B(N1390));
XOR2XL inst_blk01_cellmath__39_I877 (.Y(N1840), .A(N1392), .B(N1390));
XOR2XL inst_blk01_cellmath__39_I879 (.Y(N1842), .A(N1394), .B(N1393));
NOR2XL inst_blk01_cellmath__39_I880 (.Y(N1843), .A(N1395), .B(N1396));
XOR2XL inst_blk01_cellmath__39_I881 (.Y(N1844), .A(N1395), .B(N1396));
XOR2XL inst_blk01_cellmath__39_I883 (.Y(N1846), .A(N394), .B(N1397));
XNOR2X1 inst_blk01_cellmath__39_I885 (.Y(N2051), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[21]));
AOI2BB2X1 inst_blk01_cellmath__39_I1349 (.Y(N1849), .A0N(N1136), .A1N(N1143), .B0(N1779), .B1(N1782));
AOI2BB2X1 inst_blk01_cellmath__39_I1350 (.Y(N1851), .A0N(N1152), .A1N(N1159), .B0(N1783), .B1(N1786));
NAND2XL inst_blk01_cellmath__39_I889 (.Y(N1852), .A(N1786), .B(N1784));
AOI2BB2X1 inst_blk01_cellmath__39_I1351 (.Y(N1853), .A0N(N1168), .A1N(N1177), .B0(N1787), .B1(N1790));
NAND2XL inst_blk01_cellmath__39_I891 (.Y(N1854), .A(N1790), .B(N1788));
AOI2BB2X1 inst_blk01_cellmath__39_I1352 (.Y(N1855), .A0N(N1187), .A1N(N1198), .B0(N1791), .B1(N1794));
NAND2XL inst_blk01_cellmath__39_I893 (.Y(N1856), .A(N1794), .B(N1792));
AOI2BB2X1 inst_blk01_cellmath__39_I1353 (.Y(N1857), .A0N(N1211), .A1N(N1219), .B0(N1795), .B1(N1798));
NAND2XL inst_blk01_cellmath__39_I895 (.Y(N1858), .A(N1798), .B(N1796));
AOI2BB2X1 inst_blk01_cellmath__39_I1354 (.Y(N1859), .A0N(N1232), .A1N(N1243), .B0(N1799), .B1(N1802));
NAND2XL inst_blk01_cellmath__39_I897 (.Y(N1860), .A(N1802), .B(N1800));
AOI2BB2X1 inst_blk01_cellmath__39_I1355 (.Y(N1861), .A0N(N1255), .A1N(N1267), .B0(N1803), .B1(N1806));
NAND2XL inst_blk01_cellmath__39_I899 (.Y(N1862), .A(N1806), .B(N1804));
AOI2BB2X1 inst_blk01_cellmath__39_I1356 (.Y(N1863), .A0N(N1277), .A1N(N1286), .B0(N1807), .B1(N1810));
NAND2XL inst_blk01_cellmath__39_I901 (.Y(N1864), .A(N1810), .B(N1808));
AOI2BB2X1 inst_blk01_cellmath__39_I1357 (.Y(N1865), .A0N(N1297), .A1N(N1306), .B0(N1811), .B1(N1814));
NAND2XL inst_blk01_cellmath__39_I903 (.Y(N1866), .A(N1814), .B(N1812));
AOI2BB2X1 inst_blk01_cellmath__39_I1358 (.Y(N1867), .A0N(N1317), .A1N(N1324), .B0(N1815), .B1(N1818));
NAND2XL inst_blk01_cellmath__39_I905 (.Y(N1868), .A(N1818), .B(N1816));
AOI2BB2X1 inst_blk01_cellmath__39_I1359 (.Y(N1869), .A0N(N1335), .A1N(N1340), .B0(N1819), .B1(N1822));
NAND2XL inst_blk01_cellmath__39_I907 (.Y(N1870), .A(N1822), .B(N1820));
AOI2BB2X1 inst_blk01_cellmath__39_I1360 (.Y(N1871), .A0N(N1352), .A1N(N1348), .B0(N1823), .B1(N1826));
NAND2XL inst_blk01_cellmath__39_I909 (.Y(N1872), .A(N1826), .B(N1824));
AOI2BB2X1 inst_blk01_cellmath__39_I1361 (.Y(N1873), .A0N(N1360), .A1N(N1366), .B0(N1827), .B1(N1830));
NAND2XL inst_blk01_cellmath__39_I911 (.Y(N1874), .A(N1830), .B(N1828));
AOI2BB2X1 inst_blk01_cellmath__39_I1362 (.Y(N1875), .A0N(N1374), .A1N(N1380), .B0(N1831), .B1(N1834));
NAND2XL inst_blk01_cellmath__39_I913 (.Y(N1876), .A(N1834), .B(N1832));
AOI2BB2X1 inst_blk01_cellmath__39_I1363 (.Y(N1877), .A0N(N1388), .A1N(N1389), .B0(N1835), .B1(N1838));
NAND2XL inst_blk01_cellmath__39_I915 (.Y(N1878), .A(N1838), .B(N1836));
AOI2BB2X1 inst_blk01_cellmath__39_I1364 (.Y(N1879), .A0N(N1394), .A1N(N1393), .B0(N1839), .B1(N1842));
NAND2XL inst_blk01_cellmath__39_I917 (.Y(N1880), .A(N1842), .B(N1840));
OAI21XL inst_blk01_cellmath__39_I920 (.Y(N1883), .A0(N1852), .A1(N1849), .B0(N1851));
OAI21XL inst_blk01_cellmath__39_I922 (.Y(N1885), .A0(N1856), .A1(N1853), .B0(N1855));
NOR2XL inst_blk01_cellmath__39_I923 (.Y(N1886), .A(N1856), .B(N1854));
OAI21XL inst_blk01_cellmath__39_I924 (.Y(N1887), .A0(N1860), .A1(N1857), .B0(N1859));
NOR2XL inst_blk01_cellmath__39_I925 (.Y(N1888), .A(N1860), .B(N1858));
OAI21XL inst_blk01_cellmath__39_I926 (.Y(N1889), .A0(N1864), .A1(N1861), .B0(N1863));
NOR2XL inst_blk01_cellmath__39_I927 (.Y(N1890), .A(N1864), .B(N1862));
OAI21XL inst_blk01_cellmath__39_I928 (.Y(N1891), .A0(N1868), .A1(N1865), .B0(N1867));
NOR2XL inst_blk01_cellmath__39_I929 (.Y(N1892), .A(N1868), .B(N1866));
OAI21XL inst_blk01_cellmath__39_I930 (.Y(N1893), .A0(N1872), .A1(N1869), .B0(N1871));
NOR2XL inst_blk01_cellmath__39_I931 (.Y(N1894), .A(N1872), .B(N1870));
OAI21XL inst_blk01_cellmath__39_I932 (.Y(N1895), .A0(N1876), .A1(N1873), .B0(N1875));
NOR2XL inst_blk01_cellmath__39_I933 (.Y(N1896), .A(N1876), .B(N1874));
OAI21XL inst_blk01_cellmath__39_I934 (.Y(N1897), .A0(N1880), .A1(N1877), .B0(N1879));
NOR2XL inst_blk01_cellmath__39_I935 (.Y(N1898), .A(N1880), .B(N1878));
AOI21XL inst_blk01_cellmath__39_I936 (.Y(N1899), .A0(N1886), .A1(N1883), .B0(N1885));
AOI21XL inst_blk01_cellmath__39_I938 (.Y(N1901), .A0(N1890), .A1(N1887), .B0(N1889));
NAND2XL inst_blk01_cellmath__39_I939 (.Y(N1902), .A(N1890), .B(N1888));
AOI21XL inst_blk01_cellmath__39_I942 (.Y(N1905), .A0(N1898), .A1(N1895), .B0(N1897));
NAND2XL inst_blk01_cellmath__39_I943 (.Y(N1906), .A(N1898), .B(N1896));
OAI21XL inst_blk01_cellmath__39_I944 (.Y(N1907), .A0(N1902), .A1(N1899), .B0(N1901));
AO21XL inst_blk01_cellmath__39_I1366 (.Y(N1910), .A0(N1894), .A1(N1891), .B0(N1893));
AOI31X1 inst_blk01_cellmath__39_I1367 (.Y(N1911), .A0(N1894), .A1(N1892), .A2(N1907), .B0(N1910));
INVXL inst_blk01_cellmath__39_I950 (.Y(N1913), .A(N1888));
INVXL inst_blk01_cellmath__39_I951 (.Y(N1914), .A(N1887));
OAI21XL inst_blk01_cellmath__39_I952 (.Y(N1915), .A0(N1913), .A1(N1899), .B0(N1914));
INVXL inst_blk01_cellmath__39_I1506 (.Y(N3380), .A(N1907));
AOI21XL inst_blk01_cellmath__39_I956 (.Y(N1919), .A0(N1892), .A1(N1907), .B0(N1891));
INVXL inst_blk01_cellmath__39_I1507 (.Y(N3381), .A(N1911));
INVXL inst_blk01_cellmath__39_I960 (.Y(N1923), .A(N1896));
INVXL inst_blk01_cellmath__39_I961 (.Y(N1924), .A(N1895));
OAI21XL inst_blk01_cellmath__39_I962 (.Y(N1925), .A0(N1923), .A1(N1911), .B0(N1924));
OAI21XL inst_blk01_cellmath__39_I964 (.Y(N1927), .A0(N1906), .A1(N1911), .B0(N1905));
INVXL inst_blk01_cellmath__39_I966 (.Y(N1929), .A(N1854));
INVXL inst_blk01_cellmath__39_I967 (.Y(N1930), .A(N1853));
AOI21XL inst_blk01_cellmath__39_I968 (.Y(N1931), .A0(N1929), .A1(N1883), .B0(N1930));
INVXL inst_blk01_cellmath__39_I1508 (.Y(N3382), .A(N1899));
OAI21XL inst_blk01_cellmath__39_I972 (.Y(N1935), .A0(N1858), .A1(N1899), .B0(N1857));
INVXL inst_blk01_cellmath__39_I1509 (.Y(N3383), .A(N1915));
INVXL inst_blk01_cellmath__39_I976 (.Y(N1939), .A(N1862));
INVXL inst_blk01_cellmath__39_I977 (.Y(N1940), .A(N1861));
AOI21XL inst_blk01_cellmath__39_I978 (.Y(N1941), .A0(N1939), .A1(N1915), .B0(N1940));
INVXL inst_blk01_cellmath__39_I1510 (.Y(N3384), .A(N3380));
OAI21XL inst_blk01_cellmath__39_I982 (.Y(N1945), .A0(N1866), .A1(N3380), .B0(N1865));
INVXL inst_blk01_cellmath__39_I1511 (.Y(N3385), .A(N1919));
OAI21XL inst_blk01_cellmath__39_I986 (.Y(N1949), .A0(N1870), .A1(N1919), .B0(N1869));
INVXL inst_blk01_cellmath__39_I1512 (.Y(N3386), .A(N3381));
INVXL inst_blk01_cellmath__39_I990 (.Y(N1953), .A(N1874));
INVXL inst_blk01_cellmath__39_I991 (.Y(N1954), .A(N1873));
AOI21XL inst_blk01_cellmath__39_I992 (.Y(N1955), .A0(N1953), .A1(N3381), .B0(N1954));
INVXL inst_blk01_cellmath__39_I1513 (.Y(N3387), .A(N1925));
INVXL inst_blk01_cellmath__39_I996 (.Y(N1959), .A(N1878));
INVXL inst_blk01_cellmath__39_I997 (.Y(N1960), .A(N1877));
AOI21XL inst_blk01_cellmath__39_I998 (.Y(N1961), .A0(N1959), .A1(N1925), .B0(N1960));
INVXL inst_blk01_cellmath__39_I1514 (.Y(N3388), .A(N1927));
OAI2BB2XL inst_blk01_cellmath__39_I1368 (.Y(N1966), .A0N(N1843), .A1N(N1846), .B0(N394), .B1(N1397));
AOI31X1 inst_blk01_cellmath__39_I1369 (.Y(N1967), .A0(N1846), .A1(N1844), .A2(N1927), .B0(N1966));
INVXL inst_blk01_cellmath__39_I1006 (.Y(N1969), .A(N1784));
INVXL inst_blk01_cellmath__39_I1007 (.Y(N1970), .A(N1783));
OAI21XL inst_blk01_cellmath__39_I1008 (.Y(N1971), .A0(N1969), .A1(N1849), .B0(N1970));
AOI21XL inst_blk01_cellmath__39_I1012 (.Y(N1975), .A0(N1788), .A1(N1883), .B0(N1787));
INVXL inst_blk01_cellmath__39_I1016 (.Y(N1979), .A(N1792));
INVXL inst_blk01_cellmath__39_I1017 (.Y(N1980), .A(N1791));
OAI21XL inst_blk01_cellmath__39_I1018 (.Y(N1981), .A0(N1979), .A1(N1931), .B0(N1980));
AOI21XL inst_blk01_cellmath__39_I1022 (.Y(N1985), .A0(N1796), .A1(N3382), .B0(N1795));
AOI21XL inst_blk01_cellmath__39_I1026 (.Y(N1989), .A0(N1800), .A1(N1935), .B0(N1799));
INVXL inst_blk01_cellmath__39_I1030 (.Y(N1993), .A(N1804));
INVXL inst_blk01_cellmath__39_I1031 (.Y(N1994), .A(N1803));
OAI21XL inst_blk01_cellmath__39_I1032 (.Y(N1995), .A0(N1993), .A1(N3383), .B0(N1994));
INVXL inst_blk01_cellmath__39_I1036 (.Y(N1999), .A(N1808));
INVXL inst_blk01_cellmath__39_I1037 (.Y(N2000), .A(N1807));
OAI21XL inst_blk01_cellmath__39_I1038 (.Y(N2001), .A0(N1999), .A1(N1941), .B0(N2000));
AOI21XL inst_blk01_cellmath__39_I1042 (.Y(N2005), .A0(N1812), .A1(N3384), .B0(N1811));
AOI21XL inst_blk01_cellmath__39_I1046 (.Y(N2009), .A0(N1816), .A1(N1945), .B0(N1815));
AOI21XL inst_blk01_cellmath__39_I1050 (.Y(N2013), .A0(N1820), .A1(N3385), .B0(N1819));
AOI21XL inst_blk01_cellmath__39_I1054 (.Y(N2017), .A0(N1824), .A1(N1949), .B0(N1823));
INVXL inst_blk01_cellmath__39_I1058 (.Y(N2021), .A(N1828));
INVXL inst_blk01_cellmath__39_I1059 (.Y(N2022), .A(N1827));
OAI21XL inst_blk01_cellmath__39_I1060 (.Y(N2023), .A0(N2021), .A1(N3386), .B0(N2022));
INVXL inst_blk01_cellmath__39_I1064 (.Y(N2027), .A(N1832));
INVXL inst_blk01_cellmath__39_I1065 (.Y(N2028), .A(N1831));
OAI21XL inst_blk01_cellmath__39_I1066 (.Y(N2029), .A0(N2027), .A1(N1955), .B0(N2028));
INVXL inst_blk01_cellmath__39_I1070 (.Y(N2033), .A(N1836));
INVXL inst_blk01_cellmath__39_I1071 (.Y(N2034), .A(N1835));
OAI21XL inst_blk01_cellmath__39_I1072 (.Y(N2035), .A0(N2033), .A1(N3387), .B0(N2034));
INVXL inst_blk01_cellmath__39_I1076 (.Y(N2039), .A(N1840));
INVXL inst_blk01_cellmath__39_I1077 (.Y(N2040), .A(N1839));
OAI21XL inst_blk01_cellmath__39_I1078 (.Y(N2041), .A0(N2039), .A1(N1961), .B0(N2040));
INVXL inst_blk01_cellmath__39_I1082 (.Y(N2045), .A(N1844));
INVXL inst_blk01_cellmath__39_I1083 (.Y(N2046), .A(N1843));
OAI21XL inst_blk01_cellmath__39_I1084 (.Y(N2047), .A0(N2045), .A1(N3388), .B0(N2046));
XNOR2X1 inst_blk01_cellmath__39_I1096 (.Y(inst_blk01_cellmath__39_out0[20]), .A(N1779), .B(N1782));
XOR2XL inst_blk01_cellmath__39_I1097 (.Y(inst_blk01_cellmath__39_out0[21]), .A(N1849), .B(N1784));
XNOR2X1 inst_blk01_cellmath__39_I1098 (.Y(inst_blk01_cellmath__39_out0[22]), .A(N1971), .B(N1786));
XNOR2X1 inst_blk01_cellmath__39_I1099 (.Y(inst_blk01_cellmath__39_out0[23]), .A(N1883), .B(N1788));
XOR2XL inst_blk01_cellmath__39_I1100 (.Y(inst_blk01_cellmath__39_out0[24]), .A(N1975), .B(N1790));
XOR2XL inst_blk01_cellmath__39_I1556 (.Y(inst_blk01_cellmath__39_out0[25]), .A(N1931), .B(N1792));
XNOR2X1 inst_blk01_cellmath__39_I1102 (.Y(inst_blk01_cellmath__39_out0[26]), .A(N1981), .B(N1794));
XNOR2X1 inst_blk01_cellmath__39_I1103 (.Y(inst_blk01_cellmath__39_out0[27]), .A(N3382), .B(N1796));
XOR2XL inst_blk01_cellmath__39_I1104 (.Y(inst_blk01_cellmath__39_out0[28]), .A(N1985), .B(N1798));
XNOR2X1 inst_blk01_cellmath__39_I1105 (.Y(inst_blk01_cellmath__39_out0[29]), .A(N1935), .B(N1800));
XOR2XL inst_blk01_cellmath__39_I1106 (.Y(inst_blk01_cellmath__39_out0[30]), .A(N1989), .B(N1802));
XOR2XL inst_blk01_cellmath__39_I1557 (.Y(inst_blk01_cellmath__39_out0[31]), .A(N3383), .B(N1804));
XNOR2X1 inst_blk01_cellmath__39_I1108 (.Y(inst_blk01_cellmath__39_out0[32]), .A(N1995), .B(N1806));
XOR2XL inst_blk01_cellmath__39_I1558 (.Y(inst_blk01_cellmath__39_out0[33]), .A(N1941), .B(N1808));
XNOR2X1 inst_blk01_cellmath__39_I1110 (.Y(inst_blk01_cellmath__39_out0[34]), .A(N2001), .B(N1810));
XNOR2X1 inst_blk01_cellmath__39_I1111 (.Y(inst_blk01_cellmath__39_out0[35]), .A(N3384), .B(N1812));
XOR2XL inst_blk01_cellmath__39_I1112 (.Y(inst_blk01_cellmath__39_out0[36]), .A(N2005), .B(N1814));
XNOR2X1 inst_blk01_cellmath__39_I1113 (.Y(inst_blk01_cellmath__39_out0[37]), .A(N1945), .B(N1816));
XOR2XL inst_blk01_cellmath__39_I1114 (.Y(inst_blk01_cellmath__39_out0[38]), .A(N2009), .B(N1818));
XNOR2X1 inst_blk01_cellmath__39_I1115 (.Y(inst_blk01_cellmath__39_out0[39]), .A(N3385), .B(N1820));
XOR2XL inst_blk01_cellmath__39_I1116 (.Y(inst_blk01_cellmath__39_out0[40]), .A(N2013), .B(N1822));
XNOR2X1 inst_blk01_cellmath__39_I1117 (.Y(inst_blk01_cellmath__39_out0[41]), .A(N1949), .B(N1824));
XOR2XL inst_blk01_cellmath__39_I1118 (.Y(inst_blk01_cellmath__39_out0[42]), .A(N2017), .B(N1826));
XOR2XL inst_blk01_cellmath__39_I1559 (.Y(inst_blk01_cellmath__39_out0[43]), .A(N3386), .B(N1828));
XNOR2X1 inst_blk01_cellmath__39_I1120 (.Y(inst_blk01_cellmath__39_out0[44]), .A(N2023), .B(N1830));
XOR2XL inst_blk01_cellmath__39_I1560 (.Y(inst_blk01_cellmath__39_out0[45]), .A(N1955), .B(N1832));
XNOR2X1 inst_blk01_cellmath__39_I1122 (.Y(inst_blk01_cellmath__39_out0[46]), .A(N2029), .B(N1834));
XOR2XL inst_blk01_cellmath__39_I1561 (.Y(inst_blk01_cellmath__39_out0[47]), .A(N3387), .B(N1836));
XNOR2X1 inst_blk01_cellmath__39_I1124 (.Y(inst_blk01_cellmath__39_out0[48]), .A(N2035), .B(N1838));
XOR2XL inst_blk01_cellmath__39_I1562 (.Y(inst_blk01_cellmath__39_out0[49]), .A(N1961), .B(N1840));
XNOR2X1 inst_blk01_cellmath__39_I1126 (.Y(inst_blk01_cellmath__39_out0[50]), .A(N2041), .B(N1842));
XOR2XL inst_blk01_cellmath__39_I1563 (.Y(inst_blk01_cellmath__39_out0[51]), .A(N3388), .B(N1844));
XNOR2X1 inst_blk01_cellmath__39_I1128 (.Y(inst_blk01_cellmath__39_out0[52]), .A(N2047), .B(N1846));
XNOR2X1 inst_blk01_cellmath__39_I1129 (.Y(inst_blk01_cellmath__39_out0[53]), .A(N1967), .B(N2051));
OA22X1 inst_blk01_cellmath__39_I1371 (.Y(inst_blk01_cellmath__39_out0[55]), .A0(N2051), .A1(N1967), .B0(inst_blk01_cellmath__39_in0[22]), .B1(inst_blk01_cellmath__39_in0[21]));
INVXL inst_blk01_cellmath__39_I1523 (.Y(inst_blk01_cellmath__39_out0[54]), .A(inst_blk01_cellmath__39_out0[55]));
assign inst_blk01_cellmath__39_out0[0] = 1'B0;
assign inst_blk01_cellmath__39_out0[1] = inst_blk01_cellmath__39_in0[0];
endmodule

module cynw_cm_float_cos_inst_cellmath__42_0_bdw1114505291_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0
	); /* architecture "gate_level" */ 
output [8:0] inst_cellmath__42_0_out0;
input [7:0] inst_cellmath__42_0_in0;
wire N28,N32,N62,N71,N80,N91,N104 
	;
INVXL inst_cellmath__42_0_I5 (.Y(inst_cellmath__42_0_out0[0]), .A(inst_cellmath__42_0_in0[0]));
INVXL inst_cellmath__42_0_I6 (.Y(N28), .A(inst_cellmath__42_0_in0[1]));
INVXL inst_cellmath__42_0_I8 (.Y(N32), .A(inst_cellmath__42_0_in0[3]));
NAND2BXL inst_cellmath__42_0_I31 (.Y(N62), .AN(N28), .B(inst_cellmath__42_0_in0[2]));
NAND2XL inst_cellmath__42_0_I37 (.Y(N71), .A(N32), .B(N62));
OR2XL inst_cellmath__42_0_I45 (.Y(N80), .A(inst_cellmath__42_0_in0[4]), .B(N71));
OR2XL inst_cellmath__42_0_I55 (.Y(N91), .A(inst_cellmath__42_0_in0[5]), .B(N80));
NOR2XL inst_cellmath__42_0_I67 (.Y(N104), .A(inst_cellmath__42_0_in0[6]), .B(N91));
INVXL inst_cellmath__42_0_I99 (.Y(inst_cellmath__42_0_out0[1]), .A(N28));
XNOR2X1 inst_cellmath__42_0_I87 (.Y(inst_cellmath__42_0_out0[2]), .A(inst_cellmath__42_0_out0[1]), .B(inst_cellmath__42_0_in0[2]));
XOR2XL inst_cellmath__42_0_I106 (.Y(inst_cellmath__42_0_out0[3]), .A(N62), .B(N32));
XOR2XL inst_cellmath__42_0_I164 (.Y(inst_cellmath__42_0_out0[4]), .A(N71), .B(inst_cellmath__42_0_in0[4]));
XOR2XL inst_cellmath__42_0_I165 (.Y(inst_cellmath__42_0_out0[5]), .A(N80), .B(inst_cellmath__42_0_in0[5]));
XOR2XL inst_cellmath__42_0_I166 (.Y(inst_cellmath__42_0_out0[6]), .A(N91), .B(inst_cellmath__42_0_in0[6]));
XOR2XL inst_cellmath__42_0_I167 (.Y(inst_cellmath__42_0_out0[7]), .A(N104), .B(inst_cellmath__42_0_in0[7]));
NOR2BX1 inst_cellmath__42_0_I168 (.Y(inst_cellmath__42_0_out0[8]), .AN(inst_cellmath__42_0_in0[7]), .B(N104));
endmodule

module cynw_cm_float_cos_inst_cellmath__48_bdw1114505291_bdw (
	inst_cellmath__48_out0,
	inst_cellmath__48_in0,
	inst_cellmath__48_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__48_out0;
input [5:0] inst_cellmath__48_in0;
input [55:26] inst_cellmath__48_in1;
wire N65,N66,N67,N68,N69,N70,N71 
	,N72,N73,N74,N75,N76,N77,N78,N79 
	,N80,N81,N82,N83,N84,N85,N86,N87 
	,N88,N89,N90,N91,N92,N93,N94,N130 
	,N131,N132,N133,N134,N135,N136,N137,N138 
	,N139,N140,N141,N142,N143,N144,N145,N146 
	,N147,N148,N149,N150,N151,N152,N153,N154 
	,N155,N156,N157,N158,N160,N196,N197,N198 
	,N199,N200,N201,N202,N203,N204,N205,N206 
	,N207,N208,N209,N210,N211,N212,N213,N214 
	,N215,N216,N217,N218,N219,N220,N221,N222 
	,N224,N226,N228,N264,N265,N266,N267,N268 
	,N269,N270,N271,N272,N273,N274,N275,N276 
	,N277,N278,N279,N280,N281,N282,N283,N284 
	,N285,N286,N288,N290,N292,N294,N296,N298 
	,N300,N336,N338,N340,N342,N344,N346,N348 
	,N350,N352,N354,N356,N358,N360,N362,N364 
	,N366,N368,N370,N372,N374,N376,N378,N380 
	,N382,N384,N386,N388,N390,N392,N394,N508 
	,N510,N511,N513,N514;
INVX1 inst_cellmath__48_I384 (.Y(N508), .A(inst_cellmath__48_in0[0]));
MXI2XL inst_cellmath__48_I2 (.Y(N65), .A(inst_cellmath__48_in1[27]), .B(inst_cellmath__48_in1[26]), .S0(N508));
MXI2XL inst_cellmath__48_I3 (.Y(N66), .A(inst_cellmath__48_in1[28]), .B(inst_cellmath__48_in1[27]), .S0(N508));
MXI2XL inst_cellmath__48_I4 (.Y(N67), .A(inst_cellmath__48_in1[29]), .B(inst_cellmath__48_in1[28]), .S0(N508));
MXI2XL inst_cellmath__48_I5 (.Y(N68), .A(inst_cellmath__48_in1[30]), .B(inst_cellmath__48_in1[29]), .S0(N508));
MXI2XL inst_cellmath__48_I6 (.Y(N69), .A(inst_cellmath__48_in1[31]), .B(inst_cellmath__48_in1[30]), .S0(N508));
MXI2XL inst_cellmath__48_I7 (.Y(N70), .A(inst_cellmath__48_in1[32]), .B(inst_cellmath__48_in1[31]), .S0(N508));
MXI2XL inst_cellmath__48_I8 (.Y(N71), .A(inst_cellmath__48_in1[33]), .B(inst_cellmath__48_in1[32]), .S0(N508));
MXI2XL inst_cellmath__48_I9 (.Y(N72), .A(inst_cellmath__48_in1[34]), .B(inst_cellmath__48_in1[33]), .S0(N508));
MXI2XL inst_cellmath__48_I10 (.Y(N73), .A(inst_cellmath__48_in1[35]), .B(inst_cellmath__48_in1[34]), .S0(N508));
MXI2XL inst_cellmath__48_I11 (.Y(N74), .A(inst_cellmath__48_in1[36]), .B(inst_cellmath__48_in1[35]), .S0(N508));
MXI2XL inst_cellmath__48_I12 (.Y(N75), .A(inst_cellmath__48_in1[37]), .B(inst_cellmath__48_in1[36]), .S0(N508));
MXI2XL inst_cellmath__48_I13 (.Y(N76), .A(inst_cellmath__48_in1[38]), .B(inst_cellmath__48_in1[37]), .S0(N508));
MXI2XL inst_cellmath__48_I14 (.Y(N77), .A(inst_cellmath__48_in1[39]), .B(inst_cellmath__48_in1[38]), .S0(N508));
MXI2XL inst_cellmath__48_I15 (.Y(N78), .A(inst_cellmath__48_in1[40]), .B(inst_cellmath__48_in1[39]), .S0(N508));
MXI2XL inst_cellmath__48_I16 (.Y(N79), .A(inst_cellmath__48_in1[41]), .B(inst_cellmath__48_in1[40]), .S0(N508));
MXI2XL inst_cellmath__48_I17 (.Y(N80), .A(inst_cellmath__48_in1[42]), .B(inst_cellmath__48_in1[41]), .S0(N508));
MXI2XL inst_cellmath__48_I18 (.Y(N81), .A(inst_cellmath__48_in1[43]), .B(inst_cellmath__48_in1[42]), .S0(N508));
MXI2XL inst_cellmath__48_I19 (.Y(N82), .A(inst_cellmath__48_in1[44]), .B(inst_cellmath__48_in1[43]), .S0(N508));
MXI2XL inst_cellmath__48_I20 (.Y(N83), .A(inst_cellmath__48_in1[45]), .B(inst_cellmath__48_in1[44]), .S0(N508));
MXI2XL inst_cellmath__48_I21 (.Y(N84), .A(inst_cellmath__48_in1[46]), .B(inst_cellmath__48_in1[45]), .S0(N508));
MXI2XL inst_cellmath__48_I22 (.Y(N85), .A(inst_cellmath__48_in1[47]), .B(inst_cellmath__48_in1[46]), .S0(N508));
MXI2XL inst_cellmath__48_I23 (.Y(N86), .A(inst_cellmath__48_in1[48]), .B(inst_cellmath__48_in1[47]), .S0(N508));
MXI2XL inst_cellmath__48_I24 (.Y(N87), .A(inst_cellmath__48_in1[49]), .B(inst_cellmath__48_in1[48]), .S0(N508));
MXI2XL inst_cellmath__48_I25 (.Y(N88), .A(inst_cellmath__48_in1[50]), .B(inst_cellmath__48_in1[49]), .S0(N508));
MXI2XL inst_cellmath__48_I26 (.Y(N89), .A(inst_cellmath__48_in1[51]), .B(inst_cellmath__48_in1[50]), .S0(N508));
MXI2XL inst_cellmath__48_I27 (.Y(N90), .A(inst_cellmath__48_in1[52]), .B(inst_cellmath__48_in1[51]), .S0(N508));
MXI2XL inst_cellmath__48_I28 (.Y(N91), .A(inst_cellmath__48_in1[53]), .B(inst_cellmath__48_in1[52]), .S0(N508));
MXI2XL inst_cellmath__48_I29 (.Y(N92), .A(inst_cellmath__48_in1[54]), .B(inst_cellmath__48_in1[53]), .S0(N508));
MXI2XL inst_cellmath__48_I30 (.Y(N93), .A(inst_cellmath__48_in1[55]), .B(inst_cellmath__48_in1[54]), .S0(N508));
NAND2XL inst_cellmath__48_I31 (.Y(N94), .A(inst_cellmath__48_in1[55]), .B(N508));
BUFX2 inst_cellmath__48_I393 (.Y(N510), .A(inst_cellmath__48_in0[1]));
MXI2XL inst_cellmath__48_I66 (.Y(N130), .A(N65), .B(N67), .S0(N510));
MXI2XL inst_cellmath__48_I67 (.Y(N131), .A(N66), .B(N68), .S0(N510));
MXI2XL inst_cellmath__48_I68 (.Y(N132), .A(N67), .B(N69), .S0(N510));
MXI2XL inst_cellmath__48_I69 (.Y(N133), .A(N68), .B(N70), .S0(N510));
MXI2XL inst_cellmath__48_I70 (.Y(N134), .A(N69), .B(N71), .S0(N510));
MXI2XL inst_cellmath__48_I71 (.Y(N135), .A(N70), .B(N72), .S0(N510));
MXI2XL inst_cellmath__48_I72 (.Y(N136), .A(N71), .B(N73), .S0(N510));
MXI2XL inst_cellmath__48_I73 (.Y(N137), .A(N72), .B(N74), .S0(N510));
MXI2XL inst_cellmath__48_I74 (.Y(N138), .A(N73), .B(N75), .S0(N510));
MXI2XL inst_cellmath__48_I75 (.Y(N139), .A(N74), .B(N76), .S0(N510));
MXI2XL inst_cellmath__48_I76 (.Y(N140), .A(N75), .B(N77), .S0(N510));
MXI2XL inst_cellmath__48_I77 (.Y(N141), .A(N76), .B(N78), .S0(N510));
MXI2XL inst_cellmath__48_I78 (.Y(N142), .A(N77), .B(N79), .S0(N510));
MXI2XL inst_cellmath__48_I79 (.Y(N143), .A(N78), .B(N80), .S0(N510));
MXI2XL inst_cellmath__48_I80 (.Y(N144), .A(N79), .B(N81), .S0(N510));
MXI2XL inst_cellmath__48_I81 (.Y(N145), .A(N80), .B(N82), .S0(N510));
MXI2XL inst_cellmath__48_I82 (.Y(N146), .A(N81), .B(N83), .S0(N510));
MXI2XL inst_cellmath__48_I83 (.Y(N147), .A(N82), .B(N84), .S0(N510));
MXI2XL inst_cellmath__48_I84 (.Y(N148), .A(N83), .B(N85), .S0(N510));
MXI2XL inst_cellmath__48_I85 (.Y(N149), .A(N84), .B(N86), .S0(N510));
MXI2XL inst_cellmath__48_I86 (.Y(N150), .A(N85), .B(N87), .S0(N510));
MXI2XL inst_cellmath__48_I87 (.Y(N151), .A(N86), .B(N88), .S0(N510));
MXI2XL inst_cellmath__48_I88 (.Y(N152), .A(N87), .B(N89), .S0(N510));
MXI2XL inst_cellmath__48_I89 (.Y(N153), .A(N88), .B(N90), .S0(N510));
MXI2XL inst_cellmath__48_I90 (.Y(N154), .A(N89), .B(N91), .S0(N510));
MXI2XL inst_cellmath__48_I91 (.Y(N155), .A(N90), .B(N92), .S0(N510));
MXI2XL inst_cellmath__48_I92 (.Y(N156), .A(N91), .B(N93), .S0(N510));
MXI2XL inst_cellmath__48_I93 (.Y(N157), .A(N92), .B(N94), .S0(N510));
NOR2XL inst_cellmath__48_I94 (.Y(N158), .A(N93), .B(N510));
NOR2XL inst_cellmath__48_I95 (.Y(N160), .A(N94), .B(N510));
INVX1 inst_cellmath__48_I387 (.Y(N511), .A(inst_cellmath__48_in0[2]));
MXI2XL inst_cellmath__48_I130 (.Y(N196), .A(N134), .B(N130), .S0(N511));
MXI2XL inst_cellmath__48_I131 (.Y(N197), .A(N135), .B(N131), .S0(N511));
MXI2XL inst_cellmath__48_I132 (.Y(N198), .A(N136), .B(N132), .S0(N511));
MXI2XL inst_cellmath__48_I133 (.Y(N199), .A(N137), .B(N133), .S0(N511));
MXI2XL inst_cellmath__48_I134 (.Y(N200), .A(N138), .B(N134), .S0(N511));
MXI2XL inst_cellmath__48_I135 (.Y(N201), .A(N139), .B(N135), .S0(N511));
MXI2XL inst_cellmath__48_I136 (.Y(N202), .A(N140), .B(N136), .S0(N511));
MXI2XL inst_cellmath__48_I137 (.Y(N203), .A(N141), .B(N137), .S0(N511));
MXI2XL inst_cellmath__48_I138 (.Y(N204), .A(N142), .B(N138), .S0(N511));
MXI2XL inst_cellmath__48_I139 (.Y(N205), .A(N143), .B(N139), .S0(N511));
MXI2XL inst_cellmath__48_I140 (.Y(N206), .A(N144), .B(N140), .S0(N511));
MXI2XL inst_cellmath__48_I141 (.Y(N207), .A(N145), .B(N141), .S0(N511));
MXI2XL inst_cellmath__48_I142 (.Y(N208), .A(N146), .B(N142), .S0(N511));
MXI2XL inst_cellmath__48_I143 (.Y(N209), .A(N147), .B(N143), .S0(N511));
MXI2XL inst_cellmath__48_I144 (.Y(N210), .A(N148), .B(N144), .S0(N511));
MXI2XL inst_cellmath__48_I145 (.Y(N211), .A(N149), .B(N145), .S0(N511));
MXI2XL inst_cellmath__48_I146 (.Y(N212), .A(N150), .B(N146), .S0(N511));
MXI2XL inst_cellmath__48_I147 (.Y(N213), .A(N151), .B(N147), .S0(N511));
MXI2XL inst_cellmath__48_I148 (.Y(N214), .A(N152), .B(N148), .S0(N511));
MXI2XL inst_cellmath__48_I149 (.Y(N215), .A(N153), .B(N149), .S0(N511));
MXI2XL inst_cellmath__48_I150 (.Y(N216), .A(N154), .B(N150), .S0(N511));
MXI2XL inst_cellmath__48_I151 (.Y(N217), .A(N155), .B(N151), .S0(N511));
MXI2XL inst_cellmath__48_I152 (.Y(N218), .A(N156), .B(N152), .S0(N511));
MXI2XL inst_cellmath__48_I153 (.Y(N219), .A(N157), .B(N153), .S0(N511));
MXI2XL inst_cellmath__48_I154 (.Y(N220), .A(N158), .B(N154), .S0(N511));
MXI2XL inst_cellmath__48_I155 (.Y(N221), .A(N160), .B(N155), .S0(N511));
NAND2XL inst_cellmath__48_I156 (.Y(N222), .A(N156), .B(N511));
NAND2XL inst_cellmath__48_I157 (.Y(N224), .A(N157), .B(N511));
NAND2XL inst_cellmath__48_I158 (.Y(N226), .A(N158), .B(N511));
NAND2XL inst_cellmath__48_I159 (.Y(N228), .A(N160), .B(N511));
BUFX2 inst_cellmath__48_I394 (.Y(N513), .A(inst_cellmath__48_in0[3]));
MXI2XL inst_cellmath__48_I194 (.Y(N264), .A(N196), .B(N204), .S0(N513));
MXI2XL inst_cellmath__48_I195 (.Y(N265), .A(N197), .B(N205), .S0(N513));
MXI2XL inst_cellmath__48_I196 (.Y(N266), .A(N198), .B(N206), .S0(N513));
MXI2XL inst_cellmath__48_I197 (.Y(N267), .A(N199), .B(N207), .S0(N513));
MXI2XL inst_cellmath__48_I198 (.Y(N268), .A(N200), .B(N208), .S0(N513));
MXI2XL inst_cellmath__48_I199 (.Y(N269), .A(N201), .B(N209), .S0(N513));
MXI2XL inst_cellmath__48_I200 (.Y(N270), .A(N202), .B(N210), .S0(N513));
MXI2XL inst_cellmath__48_I201 (.Y(N271), .A(N203), .B(N211), .S0(N513));
MXI2XL inst_cellmath__48_I202 (.Y(N272), .A(N204), .B(N212), .S0(N513));
MXI2XL inst_cellmath__48_I203 (.Y(N273), .A(N205), .B(N213), .S0(N513));
MXI2XL inst_cellmath__48_I204 (.Y(N274), .A(N206), .B(N214), .S0(N513));
MXI2XL inst_cellmath__48_I205 (.Y(N275), .A(N207), .B(N215), .S0(N513));
MXI2XL inst_cellmath__48_I206 (.Y(N276), .A(N208), .B(N216), .S0(N513));
MXI2XL inst_cellmath__48_I207 (.Y(N277), .A(N209), .B(N217), .S0(N513));
MXI2XL inst_cellmath__48_I208 (.Y(N278), .A(N210), .B(N218), .S0(N513));
MXI2XL inst_cellmath__48_I209 (.Y(N279), .A(N211), .B(N219), .S0(N513));
MXI2XL inst_cellmath__48_I210 (.Y(N280), .A(N212), .B(N220), .S0(N513));
MXI2XL inst_cellmath__48_I211 (.Y(N281), .A(N213), .B(N221), .S0(N513));
MXI2XL inst_cellmath__48_I212 (.Y(N282), .A(N214), .B(N222), .S0(N513));
MXI2XL inst_cellmath__48_I213 (.Y(N283), .A(N215), .B(N224), .S0(N513));
MXI2XL inst_cellmath__48_I214 (.Y(N284), .A(N216), .B(N226), .S0(N513));
MXI2XL inst_cellmath__48_I215 (.Y(N285), .A(N217), .B(N228), .S0(N513));
NOR2XL inst_cellmath__48_I216 (.Y(N286), .A(N218), .B(N513));
NOR2XL inst_cellmath__48_I217 (.Y(N288), .A(N219), .B(N513));
NOR2XL inst_cellmath__48_I218 (.Y(N290), .A(N220), .B(N513));
NOR2XL inst_cellmath__48_I219 (.Y(N292), .A(N221), .B(N513));
NOR2XL inst_cellmath__48_I220 (.Y(N294), .A(N222), .B(N513));
NOR2XL inst_cellmath__48_I221 (.Y(N296), .A(N224), .B(N513));
NOR2XL inst_cellmath__48_I222 (.Y(N298), .A(N226), .B(N513));
NOR2XL inst_cellmath__48_I223 (.Y(N300), .A(N228), .B(N513));
INVXL inst_cellmath__48_I390 (.Y(N514), .A(inst_cellmath__48_in0[5]));
NAND2XL inst_cellmath__48_I258 (.Y(N336), .A(N264), .B(N514));
NAND2XL inst_cellmath__48_I259 (.Y(N338), .A(N265), .B(N514));
NAND2XL inst_cellmath__48_I260 (.Y(N340), .A(N266), .B(N514));
NAND2XL inst_cellmath__48_I261 (.Y(N342), .A(N267), .B(N514));
NAND2XL inst_cellmath__48_I262 (.Y(N344), .A(N268), .B(N514));
NAND2XL inst_cellmath__48_I263 (.Y(N346), .A(N269), .B(N514));
NAND2XL inst_cellmath__48_I264 (.Y(N348), .A(N270), .B(N514));
NAND2XL inst_cellmath__48_I265 (.Y(N350), .A(N271), .B(N514));
NAND2XL inst_cellmath__48_I266 (.Y(N352), .A(N272), .B(N514));
NAND2XL inst_cellmath__48_I267 (.Y(N354), .A(N273), .B(N514));
NAND2XL inst_cellmath__48_I268 (.Y(N356), .A(N274), .B(N514));
NAND2XL inst_cellmath__48_I269 (.Y(N358), .A(N275), .B(N514));
NAND2XL inst_cellmath__48_I270 (.Y(N360), .A(N276), .B(N514));
NAND2XL inst_cellmath__48_I271 (.Y(N362), .A(N277), .B(N514));
NAND2XL inst_cellmath__48_I272 (.Y(N364), .A(N278), .B(N514));
NAND2XL inst_cellmath__48_I273 (.Y(N366), .A(N279), .B(N514));
NAND2XL inst_cellmath__48_I274 (.Y(N368), .A(N280), .B(N514));
NAND2XL inst_cellmath__48_I275 (.Y(N370), .A(N281), .B(N514));
NAND2XL inst_cellmath__48_I276 (.Y(N372), .A(N282), .B(N514));
NAND2XL inst_cellmath__48_I277 (.Y(N374), .A(N283), .B(N514));
NAND2XL inst_cellmath__48_I278 (.Y(N376), .A(N284), .B(N514));
NAND2XL inst_cellmath__48_I279 (.Y(N378), .A(N285), .B(N514));
NAND2XL inst_cellmath__48_I280 (.Y(N380), .A(N286), .B(N514));
NAND2XL inst_cellmath__48_I281 (.Y(N382), .A(N288), .B(N514));
NAND2XL inst_cellmath__48_I282 (.Y(N384), .A(N290), .B(N514));
NAND2XL inst_cellmath__48_I283 (.Y(N386), .A(N292), .B(N514));
NAND2XL inst_cellmath__48_I284 (.Y(N388), .A(N294), .B(N514));
NAND2XL inst_cellmath__48_I285 (.Y(N390), .A(N296), .B(N514));
NAND2XL inst_cellmath__48_I286 (.Y(N392), .A(N298), .B(N514));
NAND2XL inst_cellmath__48_I287 (.Y(N394), .A(N300), .B(N514));
MXI2XL inst_cellmath__48_I322 (.Y(inst_cellmath__48_out0[0]), .A(N336), .B(N368), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I323 (.Y(inst_cellmath__48_out0[1]), .A(N338), .B(N370), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I324 (.Y(inst_cellmath__48_out0[2]), .A(N340), .B(N372), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I325 (.Y(inst_cellmath__48_out0[3]), .A(N342), .B(N374), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I326 (.Y(inst_cellmath__48_out0[4]), .A(N344), .B(N376), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I327 (.Y(inst_cellmath__48_out0[5]), .A(N346), .B(N378), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I328 (.Y(inst_cellmath__48_out0[6]), .A(N348), .B(N380), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I329 (.Y(inst_cellmath__48_out0[7]), .A(N350), .B(N382), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I330 (.Y(inst_cellmath__48_out0[8]), .A(N352), .B(N384), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I331 (.Y(inst_cellmath__48_out0[9]), .A(N354), .B(N386), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I332 (.Y(inst_cellmath__48_out0[10]), .A(N356), .B(N388), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I333 (.Y(inst_cellmath__48_out0[11]), .A(N358), .B(N390), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I334 (.Y(inst_cellmath__48_out0[12]), .A(N360), .B(N392), .S0(inst_cellmath__48_in0[4]));
MXI2XL inst_cellmath__48_I335 (.Y(inst_cellmath__48_out0[13]), .A(N362), .B(N394), .S0(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I336 (.Y(inst_cellmath__48_out0[14]), .A(N364), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I337 (.Y(inst_cellmath__48_out0[15]), .A(N366), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I338 (.Y(inst_cellmath__48_out0[16]), .A(N368), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I339 (.Y(inst_cellmath__48_out0[17]), .A(N370), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I340 (.Y(inst_cellmath__48_out0[18]), .A(N372), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I341 (.Y(inst_cellmath__48_out0[19]), .A(N374), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I342 (.Y(inst_cellmath__48_out0[20]), .A(N376), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I343 (.Y(inst_cellmath__48_out0[21]), .A(N378), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I344 (.Y(inst_cellmath__48_out0[22]), .A(N380), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I345 (.Y(inst_cellmath__48_out0[23]), .A(N382), .B(inst_cellmath__48_in0[4]));
NOR2XL inst_cellmath__48_I346 (.Y(inst_cellmath__48_out0[24]), .A(N384), .B(inst_cellmath__48_in0[4]));
endmodule

module cynw_cm_float_cos_inst_cellmath__58__24__bdw1114505291_bdw (
	inst_cellmath__58__24__out0,
	inst_cellmath__58__24__in0
	); /* architecture "gate_level" */ 
output [1:0] inst_cellmath__58__24__out0;
input [24:23] inst_cellmath__58__24__in0;
INVXL inst_cellmath__58__24__I13 (.Y(inst_cellmath__58__24__out0[0]), .A(inst_cellmath__58__24__in0[23]));
XNOR2X1 inst_cellmath__58__24__I16 (.Y(inst_cellmath__58__24__out0[1]), .A(inst_cellmath__58__24__in0[24]), .B(inst_cellmath__58__24__out0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__61_0_bdw1114505291_bdw (
	inst_cellmath__61_0_out0,
	inst_cellmath__61_0_in0,
	inst_cellmath__61_0_in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__61_0_out0;
input [0:0] inst_cellmath__61_0_in0;
input [22:0] inst_cellmath__61_0_in1;
wire N359;
INVXL inst_cellmath__61_0_I74 (.Y(N359), .A(inst_cellmath__61_0_in0[0]));
XNOR2X1 inst_cellmath__61_0_I27 (.Y(inst_cellmath__61_0_out0[0]), .A(inst_cellmath__61_0_in1[0]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I28 (.Y(inst_cellmath__61_0_out0[1]), .A(inst_cellmath__61_0_in1[1]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I29 (.Y(inst_cellmath__61_0_out0[2]), .A(inst_cellmath__61_0_in1[2]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I30 (.Y(inst_cellmath__61_0_out0[3]), .A(inst_cellmath__61_0_in1[3]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I31 (.Y(inst_cellmath__61_0_out0[4]), .A(inst_cellmath__61_0_in1[4]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I32 (.Y(inst_cellmath__61_0_out0[5]), .A(inst_cellmath__61_0_in1[5]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I33 (.Y(inst_cellmath__61_0_out0[6]), .A(inst_cellmath__61_0_in1[6]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I34 (.Y(inst_cellmath__61_0_out0[7]), .A(inst_cellmath__61_0_in1[7]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I35 (.Y(inst_cellmath__61_0_out0[8]), .A(inst_cellmath__61_0_in1[8]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I36 (.Y(inst_cellmath__61_0_out0[9]), .A(inst_cellmath__61_0_in1[9]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I37 (.Y(inst_cellmath__61_0_out0[10]), .A(inst_cellmath__61_0_in1[10]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I38 (.Y(inst_cellmath__61_0_out0[11]), .A(inst_cellmath__61_0_in1[11]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I39 (.Y(inst_cellmath__61_0_out0[12]), .A(inst_cellmath__61_0_in1[12]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I40 (.Y(inst_cellmath__61_0_out0[13]), .A(inst_cellmath__61_0_in1[13]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I41 (.Y(inst_cellmath__61_0_out0[14]), .A(inst_cellmath__61_0_in1[14]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I42 (.Y(inst_cellmath__61_0_out0[15]), .A(inst_cellmath__61_0_in1[15]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I43 (.Y(inst_cellmath__61_0_out0[16]), .A(inst_cellmath__61_0_in1[16]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I44 (.Y(inst_cellmath__61_0_out0[17]), .A(inst_cellmath__61_0_in1[17]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I45 (.Y(inst_cellmath__61_0_out0[18]), .A(inst_cellmath__61_0_in1[18]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I46 (.Y(inst_cellmath__61_0_out0[19]), .A(inst_cellmath__61_0_in1[19]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I47 (.Y(inst_cellmath__61_0_out0[20]), .A(inst_cellmath__61_0_in1[20]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I48 (.Y(inst_cellmath__61_0_out0[21]), .A(inst_cellmath__61_0_in1[21]), .B(N359));
XNOR2X1 inst_cellmath__61_0_I49 (.Y(inst_cellmath__61_0_out0[22]), .A(inst_cellmath__61_0_in1[22]), .B(N359));
endmodule

module cynw_cm_float_cos_inst_cellmath__195__80__2WWMM_2WWMM_bdw1114505291_bdw (
	inst_cellmath__195__80__2WWMM_2WWMM_out0,
	inst_cellmath__195__80__2WWMM_2WWMM_in0
	); /* architecture "gate_level" */ 
output [72:0] inst_cellmath__195__80__2WWMM_2WWMM_out0;
input [22:17] inst_cellmath__195__80__2WWMM_2WWMM_in0;
wire N766,N767,N771,N772,N775,N777,N778 
	,N780,N782,N787,N788,N789,N790,N791,N792 
	,N798,N799,N800,N801,N802,N803,N810,N811 
	,N825,N826,N829,N830,N832,N837,N841,N843 
	,N844,N845,N849,N852,N854,N857,N858,N859 
	,N862,N1581,N1582,N1583,N1584,N1585,N1594,N1598 
	,N1599,N1600,N1601,N1602,N1614,N1615,N1618,N1624 
	,N1625,N1626,N1628,N1638,N1640,N1643,N1645,N1648 
	,N1649,N1651,N1653,N1656,N1659,N1660,N1667,N1668 
	,N1673,N1674,N1685,N1686,N1687,N1688,N1689,N1690 
	,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698 
	,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1712 
	,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720 
	,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1736 
	,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744 
	,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752 
	,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760 
	,N1761,N1763,N2473,N2474,N2475,N2476,N2477,N2478 
	,N2480,N2481,N2482,N2483,N2484,N2487,N2493,N2494 
	,N2503,N2504,N2507,N2509,N2515,N2518,N2525,N2550 
	,N2552,N2554,N2558,N2560,N2563,N2565,N2566,N2567 
	,N2568,N2569,N3292,N3293,N3297,N3300,N3326,N3327 
	,N3329,N3331,N3333,N3334,N3335,N3336,N3339,N3340 
	,N3360,N3361,N3373,N3377,N3399,N3400,N3401,N3402 
	,N3403,N3406,N3407,N3408,N3410,N3411,N3412,N3413 
	,N3414,N3415,N3416,N3417,N3420,N3421,N3422,N3423 
	,N3424,N3426,N3431,N3432,N3434,N3437,N3438,N3439 
	,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447 
	,N3448,N3449,N3454,N3457,N3458,N3459,N3460,N3462 
	,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470 
	,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478 
	,N3479,N3480,N3482,N3484,N3485,N3486,N3487,N3492 
	,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500 
	,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508 
	,N3509,N3510,N3511,N3512,N3516,N3517,N3518,N3519 
	,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527 
	,N3528,N3529,N3530,N3531,N3532,N3534,N3542,N3543 
	,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551 
	,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559 
	,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567 
	,N3568,N3569,N3572,N4296,N4300,N4306,N4308,N4309 
	,N4310,N4311,N4312,N4334,N4335,N4354,N4358,N4363 
	,N4364,N4366,N4374,N4375,N4378,N4389,N5141,N5159 
	,N5165,N5166,N5168,N5170,N5182,N5185,N5189,N5191 
	,N5195,N5202,N5217,N5220,N5221,N5222,N5223,N5224 
	,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232 
	,N5233,N5234,N5235,N5236,N5237,N5238,N5239,N5246 
	,N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254 
	,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262 
	,N5263,N5268,N5269,N5270,N5271,N5272,N5273,N5274 
	,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282 
	,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290 
	,N5291,N5292,N5293,N5294,N5295,N6025,N6029,N6031 
	,N6032,N6034,N6035,N6036,N6086,N6094,N6108,N6815 
	,N6844,N6852,N6860,N6900,N6907,N6926,N6927,N6928 
	,N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936 
	,N6937,N6938,N6939,N6940,N6941,N6942,N6943,N6944 
	,N6955,N6956,N6957,N6958,N6959,N6960,N6961,N6962 
	,N6963,N6964,N6965,N6966,N6967,N6970,N6971,N6972 
	,N6977,N6978,N6979,N6980,N6981,N6982,N6983,N6984 
	,N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992 
	,N6993,N6994,N6995,N6996,N6997,N6998,N7001,N7003 
	,N7004,N7005,N7006,N7007,N7008,N7014,N7015,N7016 
	,N7017,N7018,N7019,N7020,N7021,N7022,N7023,N7024 
	,N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032 
	,N7033,N7034,N7039,N7040,N7041,N7042,N7043,N7044 
	,N7045,N7046,N7047,N7048,N7049,N7050,N7051,N7052 
	,N7053,N7054,N7055,N7056,N7057,N7062,N7063,N7064 
	,N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072 
	,N7073,N7074,N7075,N7076,N7077,N7078,N7079,N7080 
	,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088 
	,N7089,N7090,N7091,N7171,N7173,N7175,N7179,N7181 
	,N7183,N7187,N7191,N7193,N7195,N7197,N7199,N7201 
	,N7203,N7205,N7207,N7209,N7211,N7213,N7215,N7217 
	,N7219,N7221,N7223,N7225,N7227,N7229,N7231,N7233 
	,N7237,N7239,N7241,N7243,N7245,N7247,N7249,N7251 
	,N7253,N7255,N7257,N7291,N7301,N7340,N7375,N7395 
	,N7444,N7497,N7571,N7621,N7643,N7668,N7715,N7716 
	,N7779,N7781,N7782,N7818,N7841,N7848,N7855;
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I4721 (.Y(N7291), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I4731 (.Y(N7301), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I149 (.Y(N7171), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B(N7291));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I155 (.Y(N7173), .A(N7301), .B(N7291));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I157 (.Y(N7175), .A(N7301), .B(N7291));
AOI22X1 inst_cellmath__195__80__2WWMM_2WWMM_I5290 (.Y(N7340), .A0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7301), .B1(N7291));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I167 (.Y(N7179), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I175 (.Y(N7181), .A(N7301), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I176 (.Y(N7183), .A(N7301), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
AOI22X1 inst_cellmath__195__80__2WWMM_2WWMM_I5291 (.Y(N7375), .A0(N7291), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7301), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I181 (.Y(N7187), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I5275 (.Y(N7395), .A(N7291), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5098 (.Y(N7668), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
INVX3 inst_cellmath__195__80__2WWMM_2WWMM_I5145 (.Y(N7715), .A(N7668));
INVX3 inst_cellmath__195__80__2WWMM_2WWMM_I4874 (.Y(N7444), .A(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I445 (.Y(N766), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I446 (.Y(N767), .A0(N7444), .A1(N7183), .B0(N7171), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I447 (.Y(N7191), .A(N7444), .B(N7301));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I448 (.Y(N771), .A0(N7444), .A1(N7183), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I449 (.Y(N772), .A(N7444), .B(N7181));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I450 (.Y(N7193), .A0(N7444), .A1(N7340), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I451 (.Y(N775), .A0(N7444), .A1(N7375), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I452 (.Y(N7195), .A0(N7444), .A1(N7181), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I453 (.Y(N777), .A0(N7444), .A1(N7291), .B0(N7175), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I454 (.Y(N778), .A(N7444), .B(N7183));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I455 (.Y(N780), .A0(N7444), .A1(N7171), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I456 (.Y(N7197), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I457 (.Y(N782), .A(N7715), .B(N7301));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I458 (.Y(N7199), .A(N7444), .B(N7301));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I459 (.Y(N787), .A0(N7444), .A1(N7340), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I460 (.Y(N788), .A0(N7444), .A1(N7175), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I461 (.Y(N789), .A0(N7444), .A1(N7395), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I462 (.Y(N790), .A0(N7444), .A1(N7340), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I463 (.Y(N791), .A0(N7444), .A1(N7175), .B0(N7179), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I464 (.Y(N792), .A(N7444), .B(N7179));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I469 (.Y(N798), .A0(N7444), .A1(N7291), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I470 (.Y(N799), .A0(N7444), .A1(N7181), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I471 (.Y(N800), .A0(N7444), .A1(N7175), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I472 (.Y(N801), .A0(N7444), .A1(N7187), .B0(N7183), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I473 (.Y(N802), .A0(N7444), .A1(N7171), .B0(N7301), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I474 (.Y(N803), .A(N7444), .B(N7175));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I475 (.Y(N7201), .A0(N7444), .A1(N7173), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I476 (.Y(N7203), .A0(N7444), .A1(N7171), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I477 (.Y(N7205), .A(N7187), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I478 (.Y(N7207), .A0(N7444), .A1(N7179), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I479 (.Y(N810), .A0(N7444), .A1(N7291), .B0(N7179), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I480 (.Y(N811), .A(N7444), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I481 (.Y(N7209), .A(N7715), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I488 (.Y(N825), .A0(N7444), .A1(N7183), .B0(N7395), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I489 (.Y(N826), .A(N7444), .B(N7171));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I490 (.Y(N829), .A0(N7444), .A1(N7179), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I491 (.Y(N830), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I492 (.Y(N7211), .A0(N7444), .A1(N7173), .B0(N7179), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I493 (.Y(N832), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7183), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I494 (.Y(N7213), .A(N7444), .B(N7187));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I495 (.Y(N7215), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I496 (.Y(N837), .A0(N7444), .A1(N7375), .B0(N7291), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I498 (.Y(N841), .A(N7183), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I499 (.Y(N843), .A0(N7444), .A1(N7173), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I500 (.Y(N844), .A0(N7444), .A1(N7187), .B0(N7179), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I501 (.Y(N845), .A(N7444), .B(N7340));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I503 (.Y(N849), .A0(N7444), .A1(N7340), .B0(N7183), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I505 (.Y(N852), .A0(N7444), .A1(N7187), .B0(N7375), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I507 (.Y(N854), .A(N7444), .B(N7173));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I508 (.Y(N857), .A0(N7444), .A1(N7173), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I509 (.Y(N858), .A0(N7444), .A1(N7187), .B0(N7175), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I510 (.Y(N859), .A(N7715), .B(N7291));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I511 (.Y(N862), .A(N7715), .B(N7375));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I512 (.Y(N7217), .A(N7715), .B(N7175));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I965 (.Y(N7219), .A(N7173), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I966 (.Y(N1581), .A0(N7444), .A1(N7171), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I967 (.Y(N1582), .A0(N7444), .A1(N7171), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I968 (.Y(N1583), .A0(N7444), .A1(N7173), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I969 (.Y(N1584), .A0(N7444), .A1(N7171), .B0(N7179), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I970 (.Y(N1585), .A(N7301), .B(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I971 (.Y(N7221), .A(N7715), .B(N7171));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I973 (.Y(N7223), .A0(N7444), .A1(N7173), .B0(N7187), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I974 (.Y(N1594), .A(N7715), .B(N7183));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I975 (.Y(N7225), .A0(N7444), .A1(N7181), .B0(N7291), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I976 (.Y(N1598), .A(N7375));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I977 (.Y(N1599), .A0(N7444), .A1(N7181), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I978 (.Y(N1600), .A0(N7444), .A1(N7301), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I979 (.Y(N1601), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I980 (.Y(N1602), .A0(N7444), .A1(N7375), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I981 (.Y(N7227), .A0(N7444), .A1(N7173), .B0(N7301), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I982 (.Y(N7229), .A(N7715), .B(N7173));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I983 (.Y(N7231), .A(N7444), .B(N7187));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I987 (.Y(N1614), .A0(N7444), .A1(N7179), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I988 (.Y(N1615), .A0(N7444), .A1(N7395), .B0(N7179), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I990 (.Y(N7233), .A0(N7444), .A1(N7175), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I991 (.Y(N1618), .A0(N7444), .A1(N7171), .B0(N7173), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I4927 (.Y(N7497), .A(N7340));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I996 (.Y(N1624), .A0(N7444), .A1(N7395), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I997 (.Y(N1625), .A0(N7444), .A1(N7340), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I998 (.Y(N1626), .A0(N7444), .A1(N7395), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1000 (.Y(N1628), .A0(N7444), .A1(N7179), .B0(N7175), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1001 (.Y(N7237), .A(N7444), .B(N7179));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1006 (.Y(N1638), .A0(N7444), .A1(N7173), .B0(N7181), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1008 (.Y(N1640), .A(N7444), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1009 (.Y(N1643), .A(N7340), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1010 (.Y(N1645), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7375), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1011 (.Y(N7239), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1012 (.Y(N1648), .A0(N7444), .A1(N7395), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1013 (.Y(N1649), .A0(N7444), .A1(N7187), .B0(N7291), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1015 (.Y(N1651), .A(N7444), .B(N7173));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1016 (.Y(N1653), .A(N7444), .B(N7181));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1017 (.Y(N1656), .A(N7444), .B(N7171));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1019 (.Y(N1659), .A0(N7444), .A1(N7375), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1020 (.Y(N1660), .A0(N7444), .A1(N7175), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1025 (.Y(N1667), .A0(N7444), .A1(N7301), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1026 (.Y(N1668), .A0(N7444), .A1(N7171), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1029 (.Y(N7241), .A0(N7444), .A1(N7340), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1030 (.Y(N1673), .A0(N7444), .A1(N7395), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1031 (.Y(N1674), .A0(N7444), .A1(N7301), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5146 (.Y(N7716), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5211 (.Y(N7781), .A(N7716));
CLKINVX4 inst_cellmath__195__80__2WWMM_2WWMM_I5001 (.Y(N7571), .A(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1037 (.Y(N1685), .A0(N7571), .A1(N788), .B0(N766), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1038 (.Y(N1686), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N767), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1039 (.Y(N1687), .A0(N7571), .A1(N7219), .B0(N7191), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1040 (.Y(N1688), .A0(N7571), .A1(N1581), .B0(N771), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1041 (.Y(N1689), .A0(N7571), .A1(N1582), .B0(N772), .B1(N7781));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5209 (.Y(N7779), .A(N7716));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1042 (.Y(N1690), .A0(N7571), .A1(N1583), .B0(N7193), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1043 (.Y(N1691), .A0(N7571), .A1(N1584), .B0(N775), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1044 (.Y(N1692), .A0(N7571), .A1(N1585), .B0(N7195), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1045 (.Y(N1693), .A0(N7571), .A1(N7221), .B0(N777), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1046 (.Y(N1694), .A0(N7571), .A1(N7191), .B0(N778), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1047 (.Y(N1695), .A0(N7571), .A1(N7223), .B0(N780), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1048 (.Y(N1696), .A0(N7571), .A1(N1594), .B0(N7197), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1049 (.Y(N1697), .A0(N7571), .A1(N7225), .B0(N782), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1050 (.Y(N1698), .A0(N7571), .A1(N1598), .B0(N7199), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1051 (.Y(N1699), .A0(N7571), .A1(N1599), .B0(N787), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1052 (.Y(N1700), .A0(N7571), .A1(N1600), .B0(N788), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1053 (.Y(N1701), .A0(N7571), .A1(N1601), .B0(N789), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1054 (.Y(N1702), .A0(N7571), .A1(N1602), .B0(N790), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1055 (.Y(N1703), .A0(N7571), .A1(N7227), .B0(N791), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1056 (.Y(N1704), .A0(N7571), .A1(N7229), .B0(N792), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1057 (.Y(N1705), .A(N7779), .B(N7231));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1060 (.Y(N1712), .A0(N7571), .A1(N7217), .B0(N7195), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1061 (.Y(N1713), .A0(N7571), .A1(N1614), .B0(N798), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1062 (.Y(N1714), .A0(N7571), .A1(N1615), .B0(N799), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1063 (.Y(N1715), .A0(N7571), .A1(N7201), .B0(N800), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1064 (.Y(N1716), .A0(N7571), .A1(N7233), .B0(N801), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1065 (.Y(N1717), .A0(N7571), .A1(N1618), .B0(N802), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1066 (.Y(N1718), .A0(N7571), .A1(N7215), .B0(N803), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1067 (.Y(N1719), .A0(N7571), .A1(N7497), .B0(N7201), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1068 (.Y(N1720), .A0(N7571), .A1(N1601), .B0(N7203), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1069 (.Y(N1721), .A0(N7571), .A1(N7715), .B0(N7205), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1070 (.Y(N1722), .A0(N7571), .A1(N1624), .B0(N7207), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1071 (.Y(N1723), .A0(N7571), .A1(N1625), .B0(N810), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1072 (.Y(N1724), .A0(N7571), .A1(N1626), .B0(N811), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1073 (.Y(N1725), .A0(N7571), .A1(N7497), .B0(N7209), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1074 (.Y(N1726), .A0(N7571), .A1(N1628), .B0(N7199), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1075 (.Y(N1727), .A(N7779), .B(N7237));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1080 (.Y(N1736), .A0(N7571), .A1(N1638), .B0(N825), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1081 (.Y(N1737), .A0(N7571), .A1(N832), .B0(N826), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1082 (.Y(N1738), .A0(N7571), .A1(N1640), .B0(N829), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1083 (.Y(N1739), .A0(N7571), .A1(N1643), .B0(N830), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1084 (.Y(N1740), .A0(N7571), .A1(N1645), .B0(N7211), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1085 (.Y(N1741), .A0(N7571), .A1(N7239), .B0(N832), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1086 (.Y(N1742), .A0(N7571), .A1(N1648), .B0(N7213), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1087 (.Y(N1743), .A0(N7571), .A1(N1649), .B0(N7215), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1088 (.Y(N1744), .A0(N7571), .A1(N7223), .B0(N837), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1089 (.Y(N1745), .A0(N7571), .A1(N1651), .B0(N826), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1090 (.Y(N1746), .A0(N7571), .A1(N1653), .B0(N841), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1091 (.Y(N1747), .A0(N7571), .A1(N1656), .B0(N843), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1092 (.Y(N1748), .A0(N7571), .A1(N7233), .B0(N844), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1093 (.Y(N1749), .A0(N7571), .A1(N1659), .B0(N845), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1094 (.Y(N1750), .A0(N7571), .A1(N1660), .B0(N7193), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1095 (.Y(N1751), .A0(N7571), .A1(N1594), .B0(N849), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1096 (.Y(N1752), .A0(N7571), .A1(N1584), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1097 (.Y(N1753), .A0(N7571), .A1(N7227), .B0(N852), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1098 (.Y(N1754), .A0(N7571), .A1(N801), .B0(N7197), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1099 (.Y(N1755), .A0(N7571), .A1(N1667), .B0(N854), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1100 (.Y(N1756), .A0(N7571), .A1(N1668), .B0(N857), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1101 (.Y(N1757), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N858), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1102 (.Y(N1758), .A0(N7571), .A1(N1600), .B0(N859), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1103 (.Y(N1759), .A0(N7571), .A1(N7241), .B0(N862), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1104 (.Y(N1760), .A0(N7571), .A1(N1673), .B0(N7217), .B1(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1105 (.Y(N1761), .A(N7571), .B(N1674));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1106 (.Y(N1763), .A(N7571), .B(N7209));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1555 (.Y(N2473), .A0(N7444), .A1(N7375), .B0(N7179), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1556 (.Y(N2474), .A0(N7444), .A1(N7395), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1557 (.Y(N2475), .A0(N7444), .A1(N7187), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1558 (.Y(N2476), .A0(N7444), .A1(N7173), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1559 (.Y(N2477), .A0(N7444), .A1(N7375), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1560 (.Y(N2478), .A0(N7444), .A1(N7181), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1562 (.Y(N2480), .A0(N7444), .A1(N7173), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1563 (.Y(N2481), .A0(N7444), .A1(N7291), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1564 (.Y(N2482), .A0(N7444), .A1(N7340), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1565 (.Y(N2483), .A0(N7444), .A1(N7175), .B0(N7183), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1566 (.Y(N2484), .A(N7444), .B(N7175));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1567 (.Y(N2487), .A(N7444), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1569 (.Y(N7243), .A0(N7444), .A1(N7187), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1571 (.Y(N2493), .A0(N7444), .A1(N7291), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1572 (.Y(N2494), .A0(N7444), .A1(N7301), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1578 (.Y(N2503), .A0(N7444), .A1(N7291), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1579 (.Y(N2504), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7291), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1582 (.Y(N2507), .A(N7444), .B(N7340));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1583 (.Y(N2509), .A0(N7444), .A1(N7301), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1587 (.Y(N2515), .A0(N7444), .A1(N7375), .B0(N7181), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1589 (.Y(N2518), .A(N7444), .B(N7375));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1592 (.Y(N2525), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1605 (.Y(N2550), .A0(N7444), .A1(N7181), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1607 (.Y(N2552), .A0(N7444), .A1(N7171), .B0(N7183), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1609 (.Y(N2554), .A0(N7444), .A1(N7395), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1613 (.Y(N2558), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1614 (.Y(N7245), .A0(N7444), .A1(N7183), .B0(N7187), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1615 (.Y(N2560), .A(N7715), .B(N7181));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1616 (.Y(N2563), .A0(N7444), .A1(N7301), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(N2565), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1619 (.Y(N2566), .A0(N7444), .A1(N7301), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1620 (.Y(N2567), .A0(N7444), .A1(N7340), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1621 (.Y(N2568), .A0(N7444), .A1(N7179), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I1622 (.Y(N2569), .A0(N7444), .A1(N7291), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2074 (.Y(N3292), .A0(N7444), .A1(N7179), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2075 (.Y(N3293), .A0(N7444), .A1(N7173), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2079 (.Y(N3297), .A0(N7444), .A1(N7340), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2081 (.Y(N3300), .A0(N7444), .A1(N7340), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2096 (.Y(N3326), .A0(N7444), .A1(N7181), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2097 (.Y(N3327), .A0(N7444), .A1(N7171), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2099 (.Y(N3329), .A0(N7444), .A1(N7175), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2101 (.Y(N3331), .A0(N7444), .A1(N7183), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2102 (.Y(N7247), .A0(N7444), .A1(N7171), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2103 (.Y(N3333), .A0(N7444), .A1(N7395), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2104 (.Y(N3334), .A0(N7444), .A1(N7291), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2105 (.Y(N3335), .A0(N7444), .A1(N7183), .B0(N7179), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2106 (.Y(N3336), .A0(N7444), .A1(N7301), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2109 (.Y(N3339), .A0(N7444), .A1(N7375), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2110 (.Y(N3340), .A0(N7444), .A1(N7395), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2111 (.Y(N7249), .A0(N7444), .A1(N7187), .B0(N7173), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2122 (.Y(N3360), .A0(N7444), .A1(N7181), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2123 (.Y(N3361), .A0(N7444), .A1(N7187), .B0(N7340), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2129 (.Y(N7251), .A(N7171), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2132 (.Y(N3373), .A0(N7444), .A1(N7340), .B0(N7179), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2134 (.Y(N3377), .A(N7715), .B(N7179));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2135 (.Y(N7253), .A0(N7444), .A1(N7375), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2147 (.Y(N3399), .A0(N7571), .A1(N1615), .B0(N2473), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2148 (.Y(N3400), .A0(N7571), .A1(N3292), .B0(N2474), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2149 (.Y(N3401), .A0(N7571), .A1(N3293), .B0(N2475), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2150 (.Y(N3402), .A0(N7571), .A1(N7241), .B0(N2476), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2151 (.Y(N3403), .A(N7571), .B(N2477));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2152 (.Y(N3406), .A0(N7571), .A1(N857), .B0(N2478), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2153 (.Y(N3407), .A0(N7571), .A1(N3297), .B0(N7241), .B1(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2154 (.Y(N3408), .A(N2480), .B(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2155 (.Y(N3410), .A0(N7571), .A1(N3300), .B0(N2481), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2156 (.Y(N3411), .A0(N7571), .A1(N2481), .B0(N2482), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2157 (.Y(N3412), .A0(N7571), .A1(N7291), .B0(N2483), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2158 (.Y(N3413), .A0(N7571), .A1(N825), .B0(N2484), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2159 (.Y(N3414), .A0(N7571), .A1(N2554), .B0(N2487), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2160 (.Y(N3415), .A0(N7571), .A1(N7221), .B0(N837), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2161 (.Y(N3416), .A0(N7571), .A1(N7209), .B0(N7243), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2162 (.Y(N3417), .A(N7571), .B(N7239));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2163 (.Y(N3420), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N2493), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2164 (.Y(N3421), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N2494), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2165 (.Y(N3422), .A0(N7571), .A1(N7444), .B0(N7205), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2166 (.Y(N3423), .A0(N7571), .A1(N7444), .B0(N7715), .B1(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2167 (.Y(N3424), .A(N7571), .B(N7444));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2168 (.Y(N3426), .A(N7781), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2170 (.Y(N3431), .A0(N7571), .A1(N3326), .B0(N2503), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2171 (.Y(N3432), .A0(N7571), .A1(N3327), .B0(N2504), .B1(N7781));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2173 (.Y(N3434), .A(N7781), .B(N3329));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2174 (.Y(N3437), .A0(N7571), .A1(N1660), .B0(N2507), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2175 (.Y(N3438), .A0(N7571), .A1(N3331), .B0(N2509), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2176 (.Y(N3439), .A0(N7571), .A1(N7247), .B0(N7221), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2177 (.Y(N3440), .A0(N7571), .A1(N3333), .B0(N7197), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2178 (.Y(N3441), .A0(N7571), .A1(N3334), .B0(N1599), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2179 (.Y(N3442), .A0(N7571), .A1(N3335), .B0(N2515), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2180 (.Y(N3443), .A0(N7571), .A1(N3336), .B0(N841), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2181 (.Y(N3444), .A0(N7571), .A1(N2493), .B0(N2518), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2182 (.Y(N3445), .A0(N7571), .A1(N2525), .B0(N7237), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2183 (.Y(N3446), .A0(N7571), .A1(N3339), .B0(N2503), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2184 (.Y(N3447), .A0(N7571), .A1(N3340), .B0(N2525), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2185 (.Y(N3448), .A0(N7571), .A1(N7249), .B0(N1667), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2186 (.Y(N3449), .A0(N7571), .A1(N7219), .B0(N7213), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2189 (.Y(N3454), .A(N7779), .B(N7213));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2190 (.Y(N3457), .A0(N7571), .A1(N811), .B0(N7211), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2191 (.Y(N3458), .A0(N7571), .A1(N2484), .B0(N2507), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2192 (.Y(N3459), .A0(N7571), .A1(N788), .B0(N7715), .B1(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2193 (.Y(N3460), .A(N7571), .B(N1624));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2194 (.Y(N3462), .A0(N7571), .A1(N7197), .B0(N7199), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2195 (.Y(N3463), .A0(N7571), .A1(N3336), .B0(N782), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2196 (.Y(N3464), .A0(N7571), .A1(N3360), .B0(N7217), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2197 (.Y(N3465), .A0(N7571), .A1(N3361), .B0(N2550), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2198 (.Y(N3466), .A0(N7571), .A1(N3360), .B0(N7207), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2199 (.Y(N3467), .A0(N7571), .A1(N7203), .B0(N2552), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2200 (.Y(N3468), .A0(N7571), .A1(N3327), .B0(N7225), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2201 (.Y(N3469), .A0(N7571), .A1(N2475), .B0(N2554), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2202 (.Y(N3470), .A0(N7571), .A1(N1599), .B0(N844), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2203 (.Y(N3471), .A0(N7571), .A1(N7251), .B0(N7207), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2204 (.Y(N3472), .A0(N7571), .A1(N790), .B0(N777), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2205 (.Y(N3473), .A0(N7571), .A1(N7213), .B0(N2558), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2206 (.Y(N3474), .A0(N7571), .A1(N3373), .B0(N7245), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2207 (.Y(N3475), .A0(N7571), .A1(N782), .B0(N2560), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2208 (.Y(N3476), .A0(N7571), .A1(N3377), .B0(N2563), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2209 (.Y(N3477), .A0(N7571), .A1(N7253), .B0(N787), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2210 (.Y(N3478), .A0(N7571), .A1(N2504), .B0(N2565), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2211 (.Y(N3479), .A0(N7571), .A1(N7233), .B0(N2566), .B1(N7781));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2212 (.Y(N3480), .A(N2567), .B(N7781));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2213 (.Y(N3482), .A(N2568), .B(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2214 (.Y(N3484), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N2569), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2215 (.Y(N3485), .A0(N7571), .A1(N7497), .B0(N7193), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2216 (.Y(N3486), .A0(N7571), .A1(N7249), .B0(N7231), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2217 (.Y(N3487), .A0(N7571), .A1(N7231), .B0(N7229), .B1(N7781));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5212 (.Y(N7782), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5248 (.Y(N7818), .A(N7782));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5051 (.Y(N7621), .A(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2221 (.Y(N3492), .A0(N7621), .A1(N3399), .B0(N1685), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2222 (.Y(N3493), .A0(N7621), .A1(N3400), .B0(N1686), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2223 (.Y(N3494), .A0(N7621), .A1(N3401), .B0(N1687), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2224 (.Y(N3495), .A0(N7621), .A1(N3402), .B0(N1688), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2225 (.Y(N3496), .A0(N7621), .A1(N3403), .B0(N1689), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2226 (.Y(N3497), .A0(N7621), .A1(N3406), .B0(N1690), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2227 (.Y(N3498), .A0(N7621), .A1(N3407), .B0(N1691), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2228 (.Y(N3499), .A0(N7621), .A1(N3408), .B0(N1692), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2229 (.Y(N3500), .A0(N7621), .A1(N3410), .B0(N1693), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2230 (.Y(N3501), .A0(N7621), .A1(N3411), .B0(N1694), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2231 (.Y(N3502), .A0(N7621), .A1(N3412), .B0(N1695), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2232 (.Y(N3503), .A0(N7621), .A1(N3413), .B0(N1696), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2233 (.Y(N3504), .A0(N7621), .A1(N3414), .B0(N1697), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2234 (.Y(N3505), .A0(N7621), .A1(N3415), .B0(N1698), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2235 (.Y(N3506), .A0(N7621), .A1(N3416), .B0(N1699), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2236 (.Y(N3507), .A0(N7621), .A1(N3417), .B0(N1700), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2237 (.Y(N3508), .A0(N7621), .A1(N3420), .B0(N1701), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2238 (.Y(N3509), .A0(N7621), .A1(N3421), .B0(N1702), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2239 (.Y(N3510), .A0(N7621), .A1(N3422), .B0(N1703), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2240 (.Y(N3511), .A0(N7621), .A1(N3423), .B0(N1704), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2241 (.Y(N3512), .A0(N7621), .A1(N3424), .B0(N1705), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2244 (.Y(N3516), .A0(N7621), .A1(N3431), .B0(N1712), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2245 (.Y(N3517), .A0(N7621), .A1(N3432), .B0(N1713), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2246 (.Y(N3518), .A0(N7621), .A1(N1717), .B0(N1714), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2247 (.Y(N3519), .A0(N7621), .A1(N3434), .B0(N1715), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2248 (.Y(N3520), .A0(N7621), .A1(N3437), .B0(N1716), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2249 (.Y(N3521), .A0(N7621), .A1(N3438), .B0(N1717), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2250 (.Y(N3522), .A0(N7621), .A1(N3439), .B0(N1718), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2251 (.Y(N3523), .A0(N7621), .A1(N3440), .B0(N1719), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2252 (.Y(N3524), .A0(N7621), .A1(N3441), .B0(N1720), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2253 (.Y(N3525), .A0(N7621), .A1(N3442), .B0(N1721), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2254 (.Y(N3526), .A0(N7621), .A1(N3443), .B0(N1722), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2255 (.Y(N3527), .A0(N7621), .A1(N3444), .B0(N1723), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2256 (.Y(N3528), .A0(N7621), .A1(N3445), .B0(N1724), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2257 (.Y(N3529), .A0(N7621), .A1(N3446), .B0(N1725), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2258 (.Y(N3530), .A0(N7621), .A1(N3447), .B0(N1726), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2259 (.Y(N3531), .A0(N7621), .A1(N3448), .B0(N1727), .B1(N7818));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2260 (.Y(N3532), .A(N7621), .B(N3449));
NAND2XL hyperpropagate_3_1_A_I5294 (.Y(N7841), .A(N7571), .B(N7219));
NOR2XL hyperpropagate_3_1_A_I5295 (.Y(N3534), .A(N7818), .B(N7841));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2264 (.Y(N3542), .A0(N7621), .A1(N3457), .B0(N1736), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2265 (.Y(N3543), .A0(N7621), .A1(N3458), .B0(N1737), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2266 (.Y(N3544), .A0(N7621), .A1(N3459), .B0(N1738), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2267 (.Y(N3545), .A0(N7621), .A1(N3460), .B0(N1739), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2268 (.Y(N3546), .A0(N7621), .A1(N3462), .B0(N1740), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2269 (.Y(N3547), .A0(N7621), .A1(N3463), .B0(N1741), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2270 (.Y(N3548), .A0(N7621), .A1(N3464), .B0(N1742), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2271 (.Y(N3549), .A0(N7621), .A1(N3465), .B0(N1743), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2272 (.Y(N3550), .A0(N7621), .A1(N3466), .B0(N1744), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2273 (.Y(N3551), .A0(N7621), .A1(N3467), .B0(N1745), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2274 (.Y(N3552), .A0(N7621), .A1(N3468), .B0(N1746), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2275 (.Y(N3553), .A0(N7621), .A1(N3469), .B0(N1747), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2276 (.Y(N3554), .A0(N7621), .A1(N3470), .B0(N1748), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2277 (.Y(N3555), .A0(N7621), .A1(N3471), .B0(N1749), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2278 (.Y(N3556), .A0(N7621), .A1(N3472), .B0(N1750), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2279 (.Y(N3557), .A0(N7621), .A1(N3473), .B0(N1751), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2280 (.Y(N3558), .A0(N7621), .A1(N3474), .B0(N1752), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2281 (.Y(N3559), .A0(N7621), .A1(N3475), .B0(N1753), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2282 (.Y(N3560), .A0(N7621), .A1(N3476), .B0(N1754), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2283 (.Y(N3561), .A0(N7621), .A1(N3477), .B0(N1755), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2284 (.Y(N3562), .A0(N7621), .A1(N3478), .B0(N1756), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2285 (.Y(N3563), .A0(N7621), .A1(N3479), .B0(N1757), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2286 (.Y(N3564), .A0(N7621), .A1(N3480), .B0(N1758), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2287 (.Y(N3565), .A0(N7621), .A1(N3482), .B0(N1759), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2288 (.Y(N3566), .A0(N7621), .A1(N3484), .B0(N1760), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2289 (.Y(N3567), .A0(N7621), .A1(N3485), .B0(N1761), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2290 (.Y(N3568), .A0(N7621), .A1(N3486), .B0(N1763), .B1(N7818));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2291 (.Y(N3569), .A(N7818), .B(N3487));
NAND2XL hyperpropagate_3_1_A_I5296 (.Y(N7848), .A(N7571), .B(N7229));
NOR2XL hyperpropagate_3_1_A_I5297 (.Y(N3572), .A(N7818), .B(N7848));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2742 (.Y(N4296), .A0(N7444), .A1(N7175), .B0(N7171), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2746 (.Y(N4300), .A(N7715), .B(N7187));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2749 (.Y(N4306), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2751 (.Y(N4308), .A0(N7444), .A1(N7395), .B0(N7183), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2752 (.Y(N4309), .A(N7395));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2753 (.Y(N4310), .A0(N7444), .A1(N7179), .B0(N7183), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2754 (.Y(N4311), .A0(N7444), .A1(N7171), .B0(N7175), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2755 (.Y(N4312), .A0(N7444), .A1(N7375), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2770 (.Y(N4334), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2771 (.Y(N4335), .A0(N7444), .A1(N7187), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2784 (.Y(N4354), .A(N7715), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2786 (.Y(N4358), .A0(N7444), .A1(N7179), .B0(N7291), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2790 (.Y(N4363), .A0(N7444), .A1(N7291), .B0(N7187), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2791 (.Y(N4364), .A0(N7444), .A1(N7395), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2793 (.Y(N4366), .A(N7179), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2796 (.Y(N4374), .A0(N7444), .A1(N7179), .B0(N7181), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2797 (.Y(N4375), .A(N7444), .B(N7291));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2798 (.Y(N4378), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7171), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2801 (.Y(N7255), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7181), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I2807 (.Y(N4389), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7340), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3269 (.Y(N5141), .A(N7444), .B(N7395));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3281 (.Y(N5159), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7179), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3287 (.Y(N5165), .A(N7187));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3288 (.Y(N5166), .A0(N7444), .A1(N7340), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3290 (.Y(N5168), .A0(N7444), .A1(N7375), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3292 (.Y(N5170), .A0(N7444), .A1(N7375), .B0(N7183), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3300 (.Y(N5182), .A0(N7444), .A1(N7171), .B0(N7187), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3303 (.Y(N5185), .A(N7175));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3306 (.Y(N5189), .A0(N7444), .A1(N7183), .B0(N7375), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3308 (.Y(N5191), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7301), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3311 (.Y(N5195), .A0(N7444), .A1(N7187), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3318 (.Y(N5202), .A0(N7444), .A1(N7301), .B0(N7375), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3329 (.Y(N5217), .A(N7175), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3331 (.Y(N5220), .A0(N7571), .A1(N2568), .B0(N7197), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3332 (.Y(N5221), .A0(N7571), .A1(N1598), .B0(N862), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3333 (.Y(N5222), .A0(N7571), .A1(N7191), .B0(N7213), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3334 (.Y(N5223), .A0(N7571), .A1(N780), .B0(N4296), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3335 (.Y(N5224), .A0(N7571), .A1(N7251), .B0(N801), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3336 (.Y(N5225), .A0(N7571), .A1(N7715), .B0(N802), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3337 (.Y(N5226), .A0(N7571), .A1(N826), .B0(N7201), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3338 (.Y(N5227), .A0(N7571), .A1(N7715), .B0(N4300), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3339 (.Y(N5228), .A0(N7571), .A1(N7215), .B0(N7444), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3340 (.Y(N5229), .A0(N7571), .A1(N7243), .B0(N7253), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3341 (.Y(N5230), .A0(N7571), .A1(N843), .B0(N4306), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3342 (.Y(N5231), .A0(N7571), .A1(N7215), .B0(N2565), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3343 (.Y(N5232), .A0(N7571), .A1(N5141), .B0(N4308), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3344 (.Y(N5233), .A0(N7571), .A1(N4335), .B0(N4309), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3345 (.Y(N5234), .A0(N7571), .A1(N1643), .B0(N4310), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3346 (.Y(N5235), .A0(N7571), .A1(N7255), .B0(N4311), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3347 (.Y(N5236), .A0(N7571), .A1(N790), .B0(N4312), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3348 (.Y(N5237), .A0(N7571), .A1(N1628), .B0(N7201), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3349 (.Y(N5238), .A0(N7571), .A1(N7237), .B0(N7223), .B1(N7779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3350 (.Y(N5239), .A(N7231), .B(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3354 (.Y(N5246), .A0(N7571), .A1(N1628), .B0(N830), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3355 (.Y(N5247), .A0(N7571), .A1(N5159), .B0(N2566), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3356 (.Y(N5248), .A0(N7571), .A1(N7201), .B0(N2569), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3357 (.Y(N5249), .A0(N7571), .A1(N7249), .B0(N2518), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3358 (.Y(N5250), .A0(N7571), .A1(N7247), .B0(N771), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3359 (.Y(N5251), .A0(N7571), .A1(N7201), .B0(N7197), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3360 (.Y(N5252), .A0(N7571), .A1(N4296), .B0(N7221), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3361 (.Y(N5253), .A0(N7571), .A1(N5165), .B0(N7199), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3362 (.Y(N5254), .A0(N7571), .A1(N5166), .B0(N4334), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3363 (.Y(N5255), .A0(N7571), .A1(N3300), .B0(N4335), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3364 (.Y(N5256), .A0(N7571), .A1(N5168), .B0(N7233), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3365 (.Y(N5257), .A0(N7571), .A1(N2493), .B0(N3292), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3366 (.Y(N5258), .A0(N7571), .A1(N5170), .B0(N7291), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3367 (.Y(N5259), .A0(N7571), .A1(N791), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3368 (.Y(N5260), .A0(N7571), .A1(N7255), .B0(N7253), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3369 (.Y(N5261), .A0(N7571), .A1(N7193), .B0(N7211), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3370 (.Y(N5262), .A0(N7571), .A1(N7233), .B0(N7229), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3371 (.Y(N5263), .A0(N7571), .A1(N7217), .B0(N7231), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3374 (.Y(N5268), .A0(N7571), .A1(N5182), .B0(N7223), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3375 (.Y(N5269), .A0(N7571), .A1(N5182), .B0(N3335), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3376 (.Y(N5270), .A0(N7571), .A1(N3339), .B0(N4354), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3377 (.Y(N5271), .A0(N7571), .A1(N5185), .B0(N7203), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3378 (.Y(N5272), .A0(N7571), .A1(N2504), .B0(N4358), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3379 (.Y(N5273), .A0(N7571), .A1(N7199), .B0(N7245), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3380 (.Y(N5274), .A0(N7571), .A1(N5189), .B0(N7193), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3381 (.Y(N5275), .A0(N7571), .A1(N7195), .B0(N1651), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3382 (.Y(N5276), .A0(N7571), .A1(N5191), .B0(N4363), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3383 (.Y(N5277), .A0(N7571), .A1(N775), .B0(N4364), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3384 (.Y(N5278), .A0(N7571), .A1(N1651), .B0(N3327), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3385 (.Y(N5279), .A0(N7571), .A1(N5195), .B0(N4366), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3386 (.Y(N5280), .A0(N7571), .A1(N3293), .B0(N1640), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3387 (.Y(N5281), .A0(N7571), .A1(N7253), .B0(N1640), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3388 (.Y(N5282), .A0(N7571), .A1(N3329), .B0(N4374), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3389 (.Y(N5283), .A0(N7571), .A1(N4311), .B0(N4375), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3390 (.Y(N5284), .A0(N7571), .A1(N3339), .B0(N4378), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3391 (.Y(N5285), .A0(N7571), .A1(N7243), .B0(N7239), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3392 (.Y(N5286), .A0(N7571), .A1(N5202), .B0(N1624), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3393 (.Y(N5287), .A0(N7571), .A1(N7227), .B0(N7255), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3394 (.Y(N5288), .A0(N7571), .A1(N7245), .B0(N3340), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3395 (.Y(N5289), .A0(N7571), .A1(N1626), .B0(N4309), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3396 (.Y(N5290), .A0(N7571), .A1(N7201), .B0(N4296), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3397 (.Y(N5291), .A0(N7571), .A1(N2552), .B0(N7301), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3398 (.Y(N5292), .A0(N7571), .A1(N2515), .B0(N1601), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3399 (.Y(N5293), .A0(N7571), .A1(N1668), .B0(N4389), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3400 (.Y(N5294), .A0(N7571), .A1(N5159), .B0(N854), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3401 (.Y(N5295), .A0(N7571), .A1(N7237), .B0(N7444), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3852 (.Y(N7257), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7181), .B1(N7715));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3856 (.Y(N6025), .A(N7444), .B(N7395));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3858 (.Y(N6029), .A0(N7444), .A1(N7175), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3860 (.Y(N6031), .A0(N7444), .A1(N7291), .B0(N7183), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3861 (.Y(N6032), .A(N7181));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3863 (.Y(N6034), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7179), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3864 (.Y(N6035), .A0(N7444), .A1(N7340), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3865 (.Y(N6036), .A0(N7444), .A1(N7179), .B0(N7187), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3901 (.Y(N6086), .A(N7171));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3908 (.Y(N6094), .A(N7444), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I3918 (.Y(N6108), .A0(N7444), .A1(N7301), .B0(N7175), .B1(N7715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I4369 (.Y(N6815), .A(N7173));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4390 (.Y(N6844), .A(N7181), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4395 (.Y(N6852), .A0(N7444), .A1(N7173), .B0(N7340), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4399 (.Y(N6860), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N7340), .B1(N7715));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4424 (.Y(N6900), .A(N7395), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4428 (.Y(N6907), .A0(N7444), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N7395), .B1(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4441 (.Y(N6926), .A0(N7571), .A1(N3334), .B0(N1653), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4442 (.Y(N6927), .A0(N7571), .A1(N1638), .B0(N3292), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4443 (.Y(N6928), .A0(N7571), .A1(N6815), .B0(N5141), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4444 (.Y(N6929), .A0(N7571), .A1(N7251), .B0(N7257), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4445 (.Y(N6930), .A0(N7571), .A1(N841), .B0(N7207), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4446 (.Y(N6931), .A0(N7571), .A1(N7251), .B0(N4358), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4447 (.Y(N6932), .A0(N7571), .A1(N5170), .B0(N2560), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4448 (.Y(N6933), .A0(N7571), .A1(N2569), .B0(N6025), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4449 (.Y(N6934), .A0(N7571), .A1(N3373), .B0(N4311), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4450 (.Y(N6935), .A0(N7571), .A1(N4335), .B0(N6029), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4451 (.Y(N6936), .A0(N7571), .A1(N7227), .B0(N789), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4452 (.Y(N6937), .A0(N7571), .A1(N7241), .B0(N6031), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4453 (.Y(N6938), .A0(N7571), .A1(N6034), .B0(N6032), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4454 (.Y(N6939), .A0(N7571), .A1(N849), .B0(N5202), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4455 (.Y(N6940), .A0(N7571), .A1(N2568), .B0(N6034), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4456 (.Y(N6941), .A0(N7571), .A1(N7205), .B0(N6035), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4457 (.Y(N6942), .A0(N7571), .A1(N7444), .B0(N6036), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4458 (.Y(N6943), .A0(N7571), .A1(N7715), .B0(N7444), .B1(N7779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4459 (.Y(N6944), .A(N7571), .B(N7444));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4464 (.Y(N6955), .A0(N7571), .A1(N6844), .B0(N7247), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4465 (.Y(N6956), .A0(N7571), .A1(N803), .B0(N7245), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4466 (.Y(N6957), .A0(N7571), .A1(N4366), .B0(N7243), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4467 (.Y(N6958), .A0(N7571), .A1(N2476), .B0(N7257), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4468 (.Y(N6959), .A0(N7571), .A1(N766), .B0(N2494), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4469 (.Y(N6960), .A0(N7571), .A1(N6852), .B0(N2563), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4470 (.Y(N6961), .A0(N7571), .A1(N7251), .B0(N7201), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4471 (.Y(N6962), .A0(N7571), .A1(N7444), .B0(N4310), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4472 (.Y(N6963), .A0(N7571), .A1(N6025), .B0(N7239), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4473 (.Y(N6964), .A0(N7571), .A1(N6860), .B0(N1643), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4474 (.Y(N6965), .A0(N7571), .A1(N7257), .B0(N6031), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4475 (.Y(N6966), .A0(N7571), .A1(N7205), .B0(N7497), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4476 (.Y(N6967), .A0(N7571), .A1(N7219), .B0(N7249), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4478 (.Y(N6970), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B0(N771), .B1(N7779));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4479 (.Y(N6971), .A0(N7571), .A1(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]), .B0(N2509), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4480 (.Y(N6972), .A0(N7571), .A1(N7715), .B0(N7237), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4484 (.Y(N6977), .A0(N7571), .A1(N5185), .B0(N4308), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4485 (.Y(N6978), .A0(N7571), .A1(N6029), .B0(N7191), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4486 (.Y(N6979), .A0(N7571), .A1(N7241), .B0(N7257), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4487 (.Y(N6980), .A0(N7571), .A1(N7193), .B0(N7257), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4488 (.Y(N6981), .A0(N7571), .A1(N4358), .B0(N4364), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4489 (.Y(N6982), .A0(N7571), .A1(N1581), .B0(N2565), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4490 (.Y(N6983), .A0(N7571), .A1(N2560), .B0(N5182), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4491 (.Y(N6984), .A0(N7571), .A1(N7249), .B0(N7247), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4492 (.Y(N6985), .A0(N7571), .A1(N7225), .B0(N7203), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4493 (.Y(N6986), .A0(N7571), .A1(N4374), .B0(N6086), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4494 (.Y(N6987), .A0(N7571), .A1(N854), .B0(N7255), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4495 (.Y(N6988), .A0(N7571), .A1(N858), .B0(N7195), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4496 (.Y(N6989), .A0(N7571), .A1(N6852), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4497 (.Y(N6990), .A0(N7571), .A1(N7209), .B0(N3300), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4498 (.Y(N6991), .A0(N7571), .A1(N6900), .B0(N7253), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4499 (.Y(N6992), .A0(N7571), .A1(N7209), .B0(N7241), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4500 (.Y(N6993), .A0(N7571), .A1(N1615), .B0(N6094), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4501 (.Y(N6994), .A0(N7571), .A1(N7203), .B0(N2525), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4502 (.Y(N6995), .A0(N7571), .A1(N6907), .B0(N7225), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4503 (.Y(N6996), .A0(N7571), .A1(N7213), .B0(N3297), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4504 (.Y(N6997), .A0(N7571), .A1(N7291), .B0(N7227), .B1(N7781));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4505 (.Y(N6998), .A(N7781), .B(N7301));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4506 (.Y(N7001), .A(N7571), .B(N7715));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4507 (.Y(N7003), .A0(N7571), .A1(N2481), .B0(N7291), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4508 (.Y(N7004), .A0(N7571), .A1(N1645), .B0(N1598), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4509 (.Y(N7005), .A0(N7571), .A1(N849), .B0(N2552), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4510 (.Y(N7006), .A0(N7571), .A1(N7211), .B0(N6108), .B1(N7781));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4511 (.Y(N7007), .A0(N7571), .A1(N5217), .B0(N7199), .B1(N7781));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4512 (.Y(N7008), .A(N7571), .B(N7209));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4515 (.Y(N7014), .A0(N7621), .A1(N6926), .B0(N5220), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4516 (.Y(N7015), .A0(N7621), .A1(N6927), .B0(N5221), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4517 (.Y(N7016), .A0(N7621), .A1(N6928), .B0(N5222), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4518 (.Y(N7017), .A0(N7621), .A1(N6929), .B0(N5223), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4519 (.Y(N7018), .A0(N7621), .A1(N6930), .B0(N5224), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4520 (.Y(N7019), .A0(N7621), .A1(N6931), .B0(N5225), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4521 (.Y(N7020), .A0(N7621), .A1(N6932), .B0(N5226), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4522 (.Y(N7021), .A0(N7621), .A1(N6933), .B0(N5227), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4523 (.Y(N7022), .A0(N7621), .A1(N6934), .B0(N5228), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4524 (.Y(N7023), .A0(N7621), .A1(N6935), .B0(N5229), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4525 (.Y(N7024), .A0(N7621), .A1(N6936), .B0(N5230), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4526 (.Y(N7025), .A0(N7621), .A1(N6937), .B0(N5231), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4527 (.Y(N7026), .A0(N7621), .A1(N6938), .B0(N5232), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4528 (.Y(N7027), .A0(N7621), .A1(N6939), .B0(N5233), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4529 (.Y(N7028), .A0(N7621), .A1(N6940), .B0(N5234), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4530 (.Y(N7029), .A0(N7621), .A1(N6941), .B0(N5235), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4531 (.Y(N7030), .A0(N7621), .A1(N6942), .B0(N5236), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4532 (.Y(N7031), .A0(N7621), .A1(N6943), .B0(N5237), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4533 (.Y(N7032), .A0(N7621), .A1(N6944), .B0(N5238), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4534 (.Y(N7033), .A0(N7621), .A1(N6944), .B0(N5239), .B1(N7818));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I5278 (.Y(N7034), .A0N(N7715), .A1N(N7779), .B0(N7621));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4538 (.Y(N7039), .A0(N7621), .A1(N6955), .B0(N5246), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4539 (.Y(N7040), .A0(N7621), .A1(N6956), .B0(N5247), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4540 (.Y(N7041), .A0(N7621), .A1(N6957), .B0(N5248), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4541 (.Y(N7042), .A0(N7621), .A1(N6958), .B0(N5249), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4542 (.Y(N7043), .A0(N7621), .A1(N6959), .B0(N5250), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4543 (.Y(N7044), .A0(N7621), .A1(N6960), .B0(N5251), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4544 (.Y(N7045), .A0(N7621), .A1(N6961), .B0(N5252), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4545 (.Y(N7046), .A0(N7621), .A1(N6962), .B0(N5253), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4546 (.Y(N7047), .A0(N7621), .A1(N6963), .B0(N5254), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4547 (.Y(N7048), .A0(N7621), .A1(N6964), .B0(N5255), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4548 (.Y(N7049), .A0(N7621), .A1(N6965), .B0(N5256), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4549 (.Y(N7050), .A0(N7621), .A1(N6966), .B0(N5257), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4550 (.Y(N7051), .A0(N7621), .A1(N6967), .B0(N5258), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4551 (.Y(N7052), .A0(N7621), .A1(N5239), .B0(N5259), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4552 (.Y(N7053), .A0(N7621), .A1(N6970), .B0(N5260), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4553 (.Y(N7054), .A0(N7621), .A1(N6971), .B0(N5261), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4554 (.Y(N7055), .A0(N7621), .A1(N6972), .B0(N5262), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4555 (.Y(N7056), .A0(N7621), .A1(N7571), .B0(N5263), .B1(N7818));
NOR2XL andori2bb1_A_I5298 (.Y(N7855), .A(N7779), .B(N792));
NOR2XL andori2bb1_A_I5299 (.Y(N7057), .A(N7855), .B(N7621));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4558 (.Y(N7062), .A0(N7621), .A1(N6977), .B0(N5268), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4559 (.Y(N7063), .A0(N7621), .A1(N6978), .B0(N5269), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4560 (.Y(N7064), .A0(N7621), .A1(N6979), .B0(N5270), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4561 (.Y(N7065), .A0(N7621), .A1(N6980), .B0(N5271), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4562 (.Y(N7066), .A0(N7621), .A1(N6981), .B0(N5272), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4563 (.Y(N7067), .A0(N7621), .A1(N6982), .B0(N5273), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4564 (.Y(N7068), .A0(N7621), .A1(N6983), .B0(N5274), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4565 (.Y(N7069), .A0(N7621), .A1(N6984), .B0(N5275), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4566 (.Y(N7070), .A0(N7621), .A1(N6985), .B0(N5276), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4567 (.Y(N7071), .A0(N7621), .A1(N6986), .B0(N5277), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4568 (.Y(N7072), .A0(N7621), .A1(N6987), .B0(N5278), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4569 (.Y(N7073), .A0(N7621), .A1(N6988), .B0(N5279), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4570 (.Y(N7074), .A0(N7621), .A1(N6989), .B0(N5280), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4571 (.Y(N7075), .A0(N7621), .A1(N6990), .B0(N5281), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4572 (.Y(N7076), .A0(N7621), .A1(N6991), .B0(N5282), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4573 (.Y(N7077), .A0(N7621), .A1(N6992), .B0(N5283), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4574 (.Y(N7078), .A0(N7621), .A1(N6993), .B0(N5284), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4575 (.Y(N7079), .A0(N7621), .A1(N6994), .B0(N5285), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4576 (.Y(N7080), .A0(N7621), .A1(N6995), .B0(N5286), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4577 (.Y(N7081), .A0(N7621), .A1(N6996), .B0(N5287), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4578 (.Y(N7082), .A0(N7621), .A1(N6997), .B0(N5288), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4579 (.Y(N7083), .A0(N7621), .A1(N6998), .B0(N5289), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4580 (.Y(N7084), .A0(N7621), .A1(N7001), .B0(N5290), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4581 (.Y(N7085), .A0(N7621), .A1(N7003), .B0(N5291), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4582 (.Y(N7086), .A0(N7621), .A1(N7004), .B0(N5292), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4583 (.Y(N7087), .A0(N7621), .A1(N7005), .B0(N5293), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4584 (.Y(N7088), .A0(N7621), .A1(N7006), .B0(N5294), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4585 (.Y(N7089), .A0(N7621), .A1(N7007), .B0(N5295), .B1(N7818));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4586 (.Y(N7090), .A0(N7621), .A1(N7008), .B0(N1727), .B1(N7818));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I5280 (.Y(N7091), .A0N(N7571), .A1N(N5217), .B0(N7818));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5073 (.Y(N7643), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4589 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[0]), .A0(N7643), .A1(N7014), .B0(N3492), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4590 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[1]), .A0(N7643), .A1(N7015), .B0(N3493), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4591 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[2]), .A0(N7643), .A1(N7016), .B0(N3494), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4592 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[3]), .A0(N7643), .A1(N7017), .B0(N3495), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4593 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[4]), .A0(N7643), .A1(N7018), .B0(N3496), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4594 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[5]), .A0(N7643), .A1(N7019), .B0(N3497), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4595 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[6]), .A0(N7643), .A1(N7020), .B0(N3498), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4596 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[7]), .A0(N7643), .A1(N7021), .B0(N3499), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4597 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[8]), .A0(N7643), .A1(N7022), .B0(N3500), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4598 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[9]), .A0(N7643), .A1(N7023), .B0(N3501), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4599 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[10]), .A0(N7643), .A1(N7024), .B0(N3502), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4600 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[11]), .A0(N7643), .A1(N7025), .B0(N3503), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4601 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[12]), .A0(N7643), .A1(N7026), .B0(N3504), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4602 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[13]), .A0(N7643), .A1(N7027), .B0(N3505), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4603 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[14]), .A0(N7643), .A1(N7028), .B0(N3506), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4604 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[15]), .A0(N7643), .A1(N7029), .B0(N3507), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4605 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[16]), .A0(N7643), .A1(N7030), .B0(N3508), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4606 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[17]), .A0(N7643), .A1(N7031), .B0(N3509), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4607 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[18]), .A0(N7643), .A1(N7032), .B0(N3510), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4608 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[19]), .A0(N7643), .A1(N7033), .B0(N3511), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4609 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[20]), .A0(N7643), .A1(N7034), .B0(N3512), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I5281 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[21]), .A0N(N7621), .A1N(N3426), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4612 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[23]), .A0(N7643), .A1(N7039), .B0(N3516), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4613 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[24]), .A0(N7643), .A1(N7040), .B0(N3517), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4614 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[25]), .A0(N7643), .A1(N7041), .B0(N3518), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4615 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[26]), .A0(N7643), .A1(N7042), .B0(N3519), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4616 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[27]), .A0(N7643), .A1(N7043), .B0(N3520), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4617 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[28]), .A0(N7643), .A1(N7044), .B0(N3521), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4618 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[29]), .A0(N7643), .A1(N7045), .B0(N3522), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4619 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[30]), .A0(N7643), .A1(N7046), .B0(N3523), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4620 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[31]), .A0(N7643), .A1(N7047), .B0(N3524), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4621 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[32]), .A0(N7643), .A1(N7048), .B0(N3525), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4622 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[33]), .A0(N7643), .A1(N7049), .B0(N3526), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4623 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[34]), .A0(N7643), .A1(N7050), .B0(N3527), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4624 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[35]), .A0(N7643), .A1(N7051), .B0(N3528), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4625 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[36]), .A0(N7643), .A1(N7052), .B0(N3529), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4626 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[37]), .A0(N7643), .A1(N7053), .B0(N3530), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4627 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[38]), .A0(N7643), .A1(N7054), .B0(N3531), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4628 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[39]), .A0(N7643), .A1(N7055), .B0(N3532), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4629 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[40]), .A0(N7643), .A1(N7056), .B0(N3534), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4630 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[41]), .A0(N7643), .A1(N7057), .B0(N3534), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
OAI2BB1X1 inst_cellmath__195__80__2WWMM_2WWMM_I5282 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[42]), .A0N(N7621), .A1N(N3454), .B0(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4632 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[43]), .A0(N7643), .A1(N7062), .B0(N3542), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4633 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[44]), .A0(N7643), .A1(N7063), .B0(N3543), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4634 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[45]), .A0(N7643), .A1(N7064), .B0(N3544), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4635 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[46]), .A0(N7643), .A1(N7065), .B0(N3545), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4636 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[47]), .A0(N7643), .A1(N7066), .B0(N3546), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4637 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[48]), .A0(N7643), .A1(N7067), .B0(N3547), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4638 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[49]), .A0(N7643), .A1(N7068), .B0(N3548), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4639 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[50]), .A0(N7643), .A1(N7069), .B0(N3549), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4640 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[51]), .A0(N7643), .A1(N7070), .B0(N3550), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4641 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[52]), .A0(N7643), .A1(N7071), .B0(N3551), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4642 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[53]), .A0(N7643), .A1(N7072), .B0(N3552), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4643 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[54]), .A0(N7643), .A1(N7073), .B0(N3553), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4644 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[55]), .A0(N7643), .A1(N7074), .B0(N3554), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4645 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[56]), .A0(N7643), .A1(N7075), .B0(N3555), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4646 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[57]), .A0(N7643), .A1(N7076), .B0(N3556), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4647 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[58]), .A0(N7643), .A1(N7077), .B0(N3557), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4648 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[59]), .A0(N7643), .A1(N7078), .B0(N3558), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4649 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[60]), .A0(N7643), .A1(N7079), .B0(N3559), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4650 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[61]), .A0(N7643), .A1(N7080), .B0(N3560), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4651 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[62]), .A0(N7643), .A1(N7081), .B0(N3561), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4652 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[63]), .A0(N7643), .A1(N7082), .B0(N3562), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4653 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[64]), .A0(N7643), .A1(N7083), .B0(N3563), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4654 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[65]), .A0(N7643), .A1(N7084), .B0(N3564), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4655 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[66]), .A0(N7643), .A1(N7085), .B0(N3565), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4656 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[67]), .A0(N7643), .A1(N7086), .B0(N3566), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4657 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[68]), .A0(N7643), .A1(N7087), .B0(N3567), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4658 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[69]), .A0(N7643), .A1(N7088), .B0(N3568), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4659 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[70]), .A0(N7643), .A1(N7089), .B0(N3569), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
AOI22XL inst_cellmath__195__80__2WWMM_2WWMM_I4660 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[71]), .A0(N7643), .A1(N7090), .B0(N3572), .B1(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4661 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[72]), .A(N7643), .B(N7091));
assign inst_cellmath__195__80__2WWMM_2WWMM_out0[22] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__198_0_bdw1114505291_bdw (
	inst_cellmath__198_0_out0,
	inst_cellmath__198_0_in0,
	inst_cellmath__198_0_in1
	); /* architecture "gate_level" */ 
output [32:0] inst_cellmath__198_0_out0;
input [15:0] inst_cellmath__198_0_in0;
input [0:0] inst_cellmath__198_0_in1;
wire N102,N106,N108,N110,N112,N114,N116 
	,N118,N120,N122,N124,N126,N128,N130,N148 
	,N150,N152,N154,N156,N158,N160,N162,N164 
	,N166,N168,N170,N172,N174,N188,N192,N194 
	,N196,N198,N200,N202,N204,N206,N208,N210 
	,N212,N214,N216,N230,N234,N236,N238,N240 
	,N242,N244,N246,N248,N250,N252,N254,N256 
	,N270,N274,N276,N278,N280,N282,N284,N286 
	,N288,N290,N292,N294,N308,N312,N314,N316 
	,N318,N320,N322,N324,N326,N328,N330,N344 
	,N348,N350,N352,N354,N356,N358,N360,N362 
	,N364,N378,N382,N384,N386,N388,N390,N392 
	,N394,N396,N410,N414,N416,N418,N420,N422 
	,N424,N426,N440,N444,N446,N448,N450,N452 
	,N454,N468,N472,N474,N476,N478,N480,N494 
	,N498,N500,N502,N504,N518,N522,N524,N526 
	,N540,N544,N546,N560,N564,N578,N598,N599 
	,N600,N601,N602,N603,N604,N605,N606,N607 
	,N608,N609,N610,N611,N612,N613,N614,N615 
	,N616,N617,N618,N619,N620,N621,N622,N623 
	,N624,N625,N626,N627,N628,N629,N630,N631 
	,N632,N635,N636,N637,N638,N639,N640,N641 
	,N642,N643,N644,N645,N646,N647,N648,N649 
	,N650,N651,N652,N653,N654,N655,N656,N657 
	,N658,N659,N660,N661,N662,N663,N664,N665 
	,N666,N667,N668,N669,N670,N671,N672,N673 
	,N674,N675,N676,N677,N678,N679,N680,N681 
	,N682,N683,N684,N685,N686,N687,N688,N689 
	,N690,N691,N692,N693,N694,N695,N696,N697 
	,N698,N699,N700,N701,N702,N703,N704,N705 
	,N706,N707,N708,N709,N710,N711,N712,N713 
	,N714,N715,N716,N717,N718,N719,N720,N721 
	,N722,N723,N724,N725,N726,N727,N728,N729 
	,N730,N731,N732,N733,N734,N735,N736,N737 
	,N738,N739,N740,N741,N742,N743,N744,N745 
	,N746,N747,N748,N749,N750,N751,N752,N753 
	,N754,N755,N756,N757,N758,N759,N760,N761 
	,N762,N763,N764,N765,N766,N767,N768,N769 
	,N770,N771,N772,N773,N774,N775,N776,N777 
	,N778,N779,N780,N781,N782,N783,N784,N785 
	,N786,N787,N788,N789,N790,N791,N792,N793 
	,N794,N795,N796,N797,N798,N799,N800,N801 
	,N802,N803,N804,N805,N806,N807,N808,N809 
	,N810,N811,N812,N813,N814,N815,N816,N817 
	,N818,N819,N820,N821,N822,N823,N824,N825 
	,N826,N827,N828,N829,N830,N831,N832,N833 
	,N834,N835,N836,N837,N838,N839,N840,N841 
	,N842,N845,N855,N863,N875,N887,N903,N919 
	,N923,N924,N941,N955,N958,N961,N964,N967 
	,N970,N973,N976,N988,N990,N991,N992,N993 
	,N994,N995,N996,N997,N998,N999,N1000,N1001 
	,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009 
	,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017 
	,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025 
	,N1026,N1027,N1028,N1029,N1034,N1036,N1037,N1038 
	,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046 
	,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054 
	,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062 
	,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070 
	,N1071,N1072,N1073,N1080,N1082,N1084,N1085,N1086 
	,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094 
	,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102 
	,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110 
	,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1128 
	,N1130,N1132,N1134,N1136,N1137,N1138,N1139,N1140 
	,N1141,N1142,N1143,N1144,N1145,N1146,N1148,N1150 
	,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159 
	,N1160,N1161,N1196,N1197,N1198,N1199,N1200,N1201 
	,N1202,N1203,N1204,N1205,N1240,N1242,N1244,N1246 
	,N1248,N1257,N1260,N1263,N1266,N1269,N1272,N1275 
	,N1278,N1281,N1284,N1287,N1290,N1293,N1296,N1299 
	,N1302,N1305,N1308,N1311,N1314,N1317,N1577,N1578 
	,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586 
	,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594 
	,N1595,N1601,N1602,N1612,N1613,N1629,N1630,N1668 
	,N1669,N1670,N1671,N1672,N1673,N1674,N1675;
INVXL inst_cellmath__198_0_I952 (.Y(N1577), .A(inst_cellmath__198_0_in0[1]));
INVXL inst_cellmath__198_0_I953 (.Y(N1578), .A(inst_cellmath__198_0_in0[2]));
INVXL inst_cellmath__198_0_I954 (.Y(N1579), .A(inst_cellmath__198_0_in0[3]));
INVXL inst_cellmath__198_0_I955 (.Y(N1580), .A(inst_cellmath__198_0_in0[4]));
INVXL inst_cellmath__198_0_I956 (.Y(N1581), .A(inst_cellmath__198_0_in0[5]));
INVXL inst_cellmath__198_0_I957 (.Y(N1582), .A(inst_cellmath__198_0_in0[6]));
INVXL inst_cellmath__198_0_I958 (.Y(N1583), .A(inst_cellmath__198_0_in0[7]));
INVXL inst_cellmath__198_0_I959 (.Y(N1584), .A(inst_cellmath__198_0_in0[8]));
INVXL inst_cellmath__198_0_I960 (.Y(N1585), .A(inst_cellmath__198_0_in0[9]));
INVXL inst_cellmath__198_0_I961 (.Y(N1586), .A(inst_cellmath__198_0_in0[10]));
INVXL inst_cellmath__198_0_I962 (.Y(N1587), .A(inst_cellmath__198_0_in0[11]));
INVXL inst_cellmath__198_0_I963 (.Y(N1588), .A(inst_cellmath__198_0_in0[12]));
INVXL inst_cellmath__198_0_I964 (.Y(N1589), .A(inst_cellmath__198_0_in0[13]));
INVXL inst_cellmath__198_0_I965 (.Y(N1590), .A(inst_cellmath__198_0_in0[14]));
INVXL inst_cellmath__198_0_I966 (.Y(N1591), .A(inst_cellmath__198_0_in0[15]));
INVXL inst_cellmath__198_0_I967 (.Y(N1592), .A(inst_cellmath__198_0_in1[0]));
INVXL inst_cellmath__198_0_I968 (.Y(N1593), .A(inst_cellmath__198_0_in0[0]));
INVXL inst_cellmath__198_0_I21 (.Y(inst_cellmath__198_0_out0[0]), .A(N1593));
OR2XL inst_cellmath__198_0_I23 (.Y(N102), .A(N1593), .B(N1577));
NOR2XL inst_cellmath__198_0_I24 (.Y(N826), .A(N1593), .B(N1578));
NOR2XL inst_cellmath__198_0_I25 (.Y(N106), .A(N1593), .B(N1579));
NOR2XL inst_cellmath__198_0_I26 (.Y(N108), .A(N1593), .B(N1580));
NOR2XL inst_cellmath__198_0_I27 (.Y(N110), .A(N1593), .B(N1581));
NOR2XL inst_cellmath__198_0_I28 (.Y(N112), .A(N1593), .B(N1582));
NOR2XL inst_cellmath__198_0_I29 (.Y(N114), .A(N1593), .B(N1583));
NOR2XL inst_cellmath__198_0_I30 (.Y(N116), .A(N1593), .B(N1584));
NOR2XL inst_cellmath__198_0_I31 (.Y(N118), .A(N1593), .B(N1585));
NOR2XL inst_cellmath__198_0_I32 (.Y(N120), .A(N1593), .B(N1586));
NOR2XL inst_cellmath__198_0_I33 (.Y(N122), .A(N1593), .B(N1587));
NOR2XL inst_cellmath__198_0_I34 (.Y(N124), .A(N1593), .B(N1588));
NOR2XL inst_cellmath__198_0_I35 (.Y(N126), .A(N1593), .B(N1589));
NOR2XL inst_cellmath__198_0_I36 (.Y(N128), .A(N1593), .B(N1590));
NOR2XL inst_cellmath__198_0_I37 (.Y(N130), .A(N1593), .B(N1591));
OR2XL inst_cellmath__198_0_I38 (.Y(N598), .A(N1593), .B(N1592));
NOR2XL inst_cellmath__198_0_I45 (.Y(N148), .A(N1577), .B(N1578));
NOR2XL inst_cellmath__198_0_I46 (.Y(N150), .A(N1577), .B(N1579));
NOR2XL inst_cellmath__198_0_I47 (.Y(N152), .A(N1577), .B(N1580));
NOR2XL inst_cellmath__198_0_I48 (.Y(N154), .A(N1577), .B(N1581));
NOR2XL inst_cellmath__198_0_I49 (.Y(N156), .A(N1577), .B(N1582));
NOR2XL inst_cellmath__198_0_I50 (.Y(N158), .A(N1577), .B(N1583));
NOR2XL inst_cellmath__198_0_I51 (.Y(N160), .A(N1577), .B(N1584));
NOR2XL inst_cellmath__198_0_I52 (.Y(N162), .A(N1577), .B(N1585));
NOR2XL inst_cellmath__198_0_I53 (.Y(N164), .A(N1577), .B(N1586));
NOR2XL inst_cellmath__198_0_I54 (.Y(N166), .A(N1577), .B(N1587));
NOR2XL inst_cellmath__198_0_I55 (.Y(N168), .A(N1577), .B(N1588));
NOR2XL inst_cellmath__198_0_I56 (.Y(N170), .A(N1577), .B(N1589));
NOR2XL inst_cellmath__198_0_I57 (.Y(N172), .A(N1577), .B(N1590));
NOR2XL inst_cellmath__198_0_I58 (.Y(N174), .A(N1577), .B(N1591));
OR2XL inst_cellmath__198_0_I59 (.Y(N599), .A(N1577), .B(N1592));
INVXL inst_cellmath__198_0_I64 (.Y(N188), .A(N1578));
NOR2XL inst_cellmath__198_0_I66 (.Y(N192), .A(N1578), .B(N1579));
NOR2XL inst_cellmath__198_0_I67 (.Y(N194), .A(N1578), .B(N1580));
NOR2XL inst_cellmath__198_0_I68 (.Y(N196), .A(N1578), .B(N1581));
NOR2XL inst_cellmath__198_0_I69 (.Y(N198), .A(N1578), .B(N1582));
NOR2XL inst_cellmath__198_0_I70 (.Y(N200), .A(N1578), .B(N1583));
NOR2XL inst_cellmath__198_0_I71 (.Y(N202), .A(N1578), .B(N1584));
NOR2XL inst_cellmath__198_0_I72 (.Y(N204), .A(N1578), .B(N1585));
NOR2XL inst_cellmath__198_0_I73 (.Y(N206), .A(N1578), .B(N1586));
NOR2XL inst_cellmath__198_0_I74 (.Y(N208), .A(N1578), .B(N1587));
NOR2XL inst_cellmath__198_0_I75 (.Y(N210), .A(N1578), .B(N1588));
NOR2XL inst_cellmath__198_0_I76 (.Y(N212), .A(N1578), .B(N1589));
NOR2XL inst_cellmath__198_0_I77 (.Y(N214), .A(N1578), .B(N1590));
NOR2XL inst_cellmath__198_0_I78 (.Y(N216), .A(N1578), .B(N1591));
OR2XL inst_cellmath__198_0_I79 (.Y(N600), .A(N1578), .B(N1592));
INVXL inst_cellmath__198_0_I84 (.Y(N230), .A(N1579));
NOR2XL inst_cellmath__198_0_I86 (.Y(N234), .A(N1579), .B(N1580));
NOR2XL inst_cellmath__198_0_I87 (.Y(N236), .A(N1579), .B(N1581));
NOR2XL inst_cellmath__198_0_I88 (.Y(N238), .A(N1579), .B(N1582));
NOR2XL inst_cellmath__198_0_I89 (.Y(N240), .A(N1579), .B(N1583));
NOR2XL inst_cellmath__198_0_I90 (.Y(N242), .A(N1579), .B(N1584));
NOR2XL inst_cellmath__198_0_I91 (.Y(N244), .A(N1579), .B(N1585));
NOR2XL inst_cellmath__198_0_I92 (.Y(N246), .A(N1579), .B(N1586));
NOR2XL inst_cellmath__198_0_I93 (.Y(N248), .A(N1579), .B(N1587));
NOR2XL inst_cellmath__198_0_I94 (.Y(N250), .A(N1579), .B(N1588));
NOR2XL inst_cellmath__198_0_I95 (.Y(N252), .A(N1579), .B(N1589));
NOR2XL inst_cellmath__198_0_I96 (.Y(N254), .A(N1579), .B(N1590));
NOR2XL inst_cellmath__198_0_I97 (.Y(N256), .A(N1579), .B(N1591));
OR2XL inst_cellmath__198_0_I98 (.Y(N601), .A(N1579), .B(N1592));
INVXL inst_cellmath__198_0_I103 (.Y(N270), .A(N1580));
NOR2XL inst_cellmath__198_0_I105 (.Y(N274), .A(N1580), .B(N1581));
NOR2XL inst_cellmath__198_0_I106 (.Y(N276), .A(N1580), .B(N1582));
NOR2XL inst_cellmath__198_0_I107 (.Y(N278), .A(N1580), .B(N1583));
NOR2XL inst_cellmath__198_0_I108 (.Y(N280), .A(N1580), .B(N1584));
NOR2XL inst_cellmath__198_0_I109 (.Y(N282), .A(N1580), .B(N1585));
NOR2XL inst_cellmath__198_0_I110 (.Y(N284), .A(N1580), .B(N1586));
NOR2XL inst_cellmath__198_0_I111 (.Y(N286), .A(N1580), .B(N1587));
NOR2XL inst_cellmath__198_0_I112 (.Y(N288), .A(N1580), .B(N1588));
NOR2XL inst_cellmath__198_0_I113 (.Y(N290), .A(N1580), .B(N1589));
NOR2XL inst_cellmath__198_0_I114 (.Y(N292), .A(N1580), .B(N1590));
NOR2XL inst_cellmath__198_0_I115 (.Y(N294), .A(N1580), .B(N1591));
OR2XL inst_cellmath__198_0_I116 (.Y(N602), .A(N1580), .B(N1592));
INVXL inst_cellmath__198_0_I121 (.Y(N308), .A(N1581));
NOR2XL inst_cellmath__198_0_I123 (.Y(N312), .A(N1581), .B(N1582));
NOR2XL inst_cellmath__198_0_I124 (.Y(N314), .A(N1581), .B(N1583));
NOR2XL inst_cellmath__198_0_I125 (.Y(N316), .A(N1581), .B(N1584));
NOR2XL inst_cellmath__198_0_I126 (.Y(N318), .A(N1581), .B(N1585));
NOR2XL inst_cellmath__198_0_I127 (.Y(N320), .A(N1581), .B(N1586));
NOR2XL inst_cellmath__198_0_I128 (.Y(N322), .A(N1581), .B(N1587));
NOR2XL inst_cellmath__198_0_I129 (.Y(N324), .A(N1581), .B(N1588));
NOR2XL inst_cellmath__198_0_I130 (.Y(N326), .A(N1581), .B(N1589));
NOR2XL inst_cellmath__198_0_I131 (.Y(N328), .A(N1581), .B(N1590));
NOR2XL inst_cellmath__198_0_I132 (.Y(N330), .A(N1581), .B(N1591));
OR2XL inst_cellmath__198_0_I133 (.Y(N603), .A(N1581), .B(N1592));
INVXL inst_cellmath__198_0_I138 (.Y(N344), .A(N1582));
NOR2XL inst_cellmath__198_0_I140 (.Y(N348), .A(N1582), .B(N1583));
NOR2XL inst_cellmath__198_0_I141 (.Y(N350), .A(N1582), .B(N1584));
NOR2XL inst_cellmath__198_0_I142 (.Y(N352), .A(N1582), .B(N1585));
NOR2XL inst_cellmath__198_0_I143 (.Y(N354), .A(N1582), .B(N1586));
NOR2XL inst_cellmath__198_0_I144 (.Y(N356), .A(N1582), .B(N1587));
NOR2XL inst_cellmath__198_0_I145 (.Y(N358), .A(N1582), .B(N1588));
NOR2XL inst_cellmath__198_0_I146 (.Y(N360), .A(N1582), .B(N1589));
NOR2XL inst_cellmath__198_0_I147 (.Y(N362), .A(N1582), .B(N1590));
NOR2XL inst_cellmath__198_0_I148 (.Y(N364), .A(N1582), .B(N1591));
OR2XL inst_cellmath__198_0_I149 (.Y(N604), .A(N1582), .B(N1592));
INVXL inst_cellmath__198_0_I154 (.Y(N378), .A(N1583));
NOR2XL inst_cellmath__198_0_I156 (.Y(N382), .A(N1583), .B(N1584));
NOR2XL inst_cellmath__198_0_I157 (.Y(N384), .A(N1583), .B(N1585));
NOR2XL inst_cellmath__198_0_I158 (.Y(N386), .A(N1583), .B(N1586));
NOR2XL inst_cellmath__198_0_I159 (.Y(N388), .A(N1583), .B(N1587));
NOR2XL inst_cellmath__198_0_I160 (.Y(N390), .A(N1583), .B(N1588));
NOR2XL inst_cellmath__198_0_I161 (.Y(N392), .A(N1583), .B(N1589));
NOR2XL inst_cellmath__198_0_I162 (.Y(N394), .A(N1583), .B(N1590));
NOR2XL inst_cellmath__198_0_I163 (.Y(N396), .A(N1583), .B(N1591));
OR2XL inst_cellmath__198_0_I164 (.Y(N605), .A(N1583), .B(N1592));
INVXL inst_cellmath__198_0_I169 (.Y(N410), .A(N1584));
NOR2XL inst_cellmath__198_0_I171 (.Y(N414), .A(N1584), .B(N1585));
NOR2XL inst_cellmath__198_0_I172 (.Y(N416), .A(N1584), .B(N1586));
NOR2XL inst_cellmath__198_0_I173 (.Y(N418), .A(N1584), .B(N1587));
NOR2XL inst_cellmath__198_0_I174 (.Y(N420), .A(N1584), .B(N1588));
NOR2XL inst_cellmath__198_0_I175 (.Y(N422), .A(N1584), .B(N1589));
NOR2XL inst_cellmath__198_0_I176 (.Y(N424), .A(N1584), .B(N1590));
NOR2XL inst_cellmath__198_0_I177 (.Y(N426), .A(N1584), .B(N1591));
OR2XL inst_cellmath__198_0_I178 (.Y(N606), .A(N1584), .B(N1592));
INVXL inst_cellmath__198_0_I183 (.Y(N440), .A(N1585));
NOR2XL inst_cellmath__198_0_I185 (.Y(N444), .A(N1585), .B(N1586));
NOR2XL inst_cellmath__198_0_I186 (.Y(N446), .A(N1585), .B(N1587));
NOR2XL inst_cellmath__198_0_I187 (.Y(N448), .A(N1585), .B(N1588));
NOR2XL inst_cellmath__198_0_I188 (.Y(N450), .A(N1585), .B(N1589));
NOR2XL inst_cellmath__198_0_I189 (.Y(N452), .A(N1585), .B(N1590));
NOR2XL inst_cellmath__198_0_I190 (.Y(N454), .A(N1585), .B(N1591));
OR2XL inst_cellmath__198_0_I191 (.Y(N607), .A(N1585), .B(N1592));
INVXL inst_cellmath__198_0_I196 (.Y(N468), .A(N1586));
NOR2XL inst_cellmath__198_0_I198 (.Y(N472), .A(N1586), .B(N1587));
NOR2XL inst_cellmath__198_0_I199 (.Y(N474), .A(N1586), .B(N1588));
NOR2XL inst_cellmath__198_0_I200 (.Y(N476), .A(N1586), .B(N1589));
NOR2XL inst_cellmath__198_0_I201 (.Y(N478), .A(N1586), .B(N1590));
NOR2XL inst_cellmath__198_0_I202 (.Y(N480), .A(N1586), .B(N1591));
OR2XL inst_cellmath__198_0_I203 (.Y(N608), .A(N1586), .B(N1592));
INVXL inst_cellmath__198_0_I208 (.Y(N494), .A(N1587));
NOR2XL inst_cellmath__198_0_I210 (.Y(N498), .A(N1587), .B(N1588));
NOR2XL inst_cellmath__198_0_I211 (.Y(N500), .A(N1587), .B(N1589));
NOR2XL inst_cellmath__198_0_I212 (.Y(N502), .A(N1587), .B(N1590));
NOR2XL inst_cellmath__198_0_I213 (.Y(N504), .A(N1587), .B(N1591));
OR2XL inst_cellmath__198_0_I214 (.Y(N609), .A(N1587), .B(N1592));
INVXL inst_cellmath__198_0_I219 (.Y(N518), .A(N1588));
NOR2XL inst_cellmath__198_0_I221 (.Y(N522), .A(N1588), .B(N1589));
NOR2XL inst_cellmath__198_0_I222 (.Y(N524), .A(N1588), .B(N1590));
NOR2XL inst_cellmath__198_0_I223 (.Y(N526), .A(N1588), .B(N1591));
OR2XL inst_cellmath__198_0_I224 (.Y(N610), .A(N1588), .B(N1592));
INVXL inst_cellmath__198_0_I229 (.Y(N540), .A(N1589));
NOR2XL inst_cellmath__198_0_I231 (.Y(N544), .A(N1589), .B(N1590));
NOR2XL inst_cellmath__198_0_I232 (.Y(N546), .A(N1589), .B(N1591));
OR2XL inst_cellmath__198_0_I233 (.Y(N611), .A(N1589), .B(N1592));
INVXL inst_cellmath__198_0_I238 (.Y(N560), .A(N1590));
NOR2XL inst_cellmath__198_0_I240 (.Y(N564), .A(N1590), .B(N1591));
OR2XL inst_cellmath__198_0_I241 (.Y(N612), .A(N1590), .B(N1592));
INVXL inst_cellmath__198_0_I246 (.Y(N578), .A(N1591));
ADDHX1 inst_cellmath__198_0_I269 (.CO(N614), .S(N613), .A(N122), .B(N312));
ADDHX1 inst_cellmath__198_0_I270 (.CO(N616), .S(N615), .A(N166), .B(N314));
ADDFX1 inst_cellmath__198_0_I271 (.CO(N618), .S(N617), .A(N126), .B(N378), .CI(N316));
ADDHX1 inst_cellmath__198_0_I272 (.CO(N620), .S(N619), .A(N246), .B(N168));
ADDFX1 inst_cellmath__198_0_I273 (.CO(N622), .S(N621), .A(N318), .B(N170), .CI(N248));
ADDHX1 inst_cellmath__198_0_I274 (.CO(N624), .S(N623), .A(N128), .B(N350));
ADDFX1 inst_cellmath__198_0_I275 (.CO(N626), .S(N625), .A(N410), .B(N130), .CI(N382));
ADDFX1 inst_cellmath__198_0_I276 (.CO(N628), .S(N627), .A(N250), .B(N320), .CI(N172));
ADDHX1 inst_cellmath__198_0_I277 (.CO(N630), .S(N629), .A(N352), .B(N286));
XNOR2X1 hap1_A_I923 (.Y(N631), .A(N174), .B(N384));
OR2XL hap1_A_I924 (.Y(N632), .A(N174), .B(N384));
ADDFX1 inst_cellmath__198_0_I279 (.CO(N636), .S(N635), .A(N252), .B(N322), .CI(N598));
ADDFX1 inst_cellmath__198_0_I280 (.CO(N638), .S(N637), .A(N288), .B(N354), .CI(N214));
ADDFX1 inst_cellmath__198_0_I281 (.CO(N640), .S(N639), .A(N599), .B(N440), .CI(N386));
ADDFX1 inst_cellmath__198_0_I282 (.CO(N642), .S(N641), .A(N254), .B(N324), .CI(N414));
ADDFX1 inst_cellmath__198_0_I283 (.CO(N644), .S(N643), .A(N290), .B(N356), .CI(N216));
ADDFX1 inst_cellmath__198_0_I284 (.CO(N646), .S(N645), .A(N326), .B(N388), .CI(N256));
ADDFX1 inst_cellmath__198_0_I285 (.CO(N648), .S(N647), .A(N358), .B(N416), .CI(N292));
ADDFX1 inst_cellmath__198_0_I286 (.CO(N650), .S(N649), .A(N601), .B(N468), .CI(N444));
ADDFX1 inst_cellmath__198_0_I287 (.CO(N652), .S(N651), .A(N328), .B(N390), .CI(N418));
ADDFX1 inst_cellmath__198_0_I288 (.CO(N654), .S(N653), .A(N392), .B(N446), .CI(N330));
ADDFX1 inst_cellmath__198_0_I289 (.CO(N656), .S(N655), .A(N603), .B(N494), .CI(N448));
ADDHX1 inst_cellmath__198_0_I290 (.CO(N658), .S(N657), .A(N114), .B(N234));
ADDHX1 inst_cellmath__198_0_I291 (.CO(N660), .S(N659), .A(N158), .B(N236));
ADDFX1 inst_cellmath__198_0_I292 (.CO(N662), .S(N661), .A(N118), .B(N308), .CI(N238));
ADDHX1 inst_cellmath__198_0_I293 (.CO(N664), .S(N663), .A(N160), .B(N274));
ADDFX1 inst_cellmath__198_0_I294 (.CO(N666), .S(N665), .A(N240), .B(N162), .CI(N120));
ADDHX1 inst_cellmath__198_0_I295 (.CO(N668), .S(N667), .A(N276), .B(N202));
ADDFX1 inst_cellmath__198_0_I296 (.CO(N670), .S(N669), .A(N242), .B(N344), .CI(N164));
ADDFX1 inst_cellmath__198_0_I297 (.CO(N672), .S(N671), .A(N204), .B(N278), .CI(N613));
ADDFX1 inst_cellmath__198_0_I298 (.CO(N674), .S(N673), .A(N124), .B(N244), .CI(N280));
ADDFX1 inst_cellmath__198_0_I299 (.CO(N676), .S(N675), .A(N614), .B(N206), .CI(N615));
ADDFX1 inst_cellmath__198_0_I300 (.CO(N678), .S(N677), .A(N282), .B(N348), .CI(N208));
ADDFX1 inst_cellmath__198_0_I301 (.CO(N680), .S(N679), .A(N619), .B(N616), .CI(N617));
ADDFX1 inst_cellmath__198_0_I302 (.CO(N682), .S(N681), .A(N210), .B(N284), .CI(N620));
ADDFX1 inst_cellmath__198_0_I303 (.CO(N684), .S(N683), .A(N623), .B(N618), .CI(N621));
ADDFX1 inst_cellmath__198_0_I304 (.CO(N686), .S(N685), .A(N624), .B(N212), .CI(N622));
ADDFX1 inst_cellmath__198_0_I305 (.CO(N688), .S(N687), .A(N625), .B(N629), .CI(N627));
ADDFX1 inst_cellmath__198_0_I306 (.CO(N690), .S(N689), .A(N631), .B(N630), .CI(N626));
ADDFX1 inst_cellmath__198_0_I307 (.CO(N692), .S(N691), .A(N635), .B(N628), .CI(N637));
ADDFX1 inst_cellmath__198_0_I308 (.CO(N694), .S(N693), .A(N636), .B(N632), .CI(N638));
ADDFX1 inst_cellmath__198_0_I309 (.CO(N696), .S(N695), .A(N641), .B(N639), .CI(N643));
ADDFX1 inst_cellmath__198_0_I310 (.CO(N698), .S(N697), .A(N640), .B(N600), .CI(N642));
ADDFX1 inst_cellmath__198_0_I311 (.CO(N700), .S(N699), .A(N645), .B(N644), .CI(N647));
ADDFX1 inst_cellmath__198_0_I312 (.CO(N702), .S(N701), .A(N294), .B(N360), .CI(N646));
ADDFX1 inst_cellmath__198_0_I313 (.CO(N704), .S(N703), .A(N649), .B(N648), .CI(N651));
ADDFX1 inst_cellmath__198_0_I314 (.CO(N706), .S(N705), .A(N362), .B(N420), .CI(N602));
ADDFX1 inst_cellmath__198_0_I315 (.CO(N708), .S(N707), .A(N652), .B(N650), .CI(N653));
ADDFX1 inst_cellmath__198_0_I316 (.CO(N710), .S(N709), .A(N472), .B(N394), .CI(N422));
ADDFX1 inst_cellmath__198_0_I317 (.CO(N712), .S(N711), .A(N654), .B(N364), .CI(N655));
ADDFX1 inst_cellmath__198_0_I318 (.CO(N714), .S(N713), .A(N396), .B(N450), .CI(N474));
ADDFX1 inst_cellmath__198_0_I319 (.CO(N716), .S(N715), .A(N604), .B(N424), .CI(N656));
ADDFX1 inst_cellmath__198_0_I320 (.CO(N718), .S(N717), .A(N605), .B(N518), .CI(N498));
ADDFX1 inst_cellmath__198_0_I321 (.CO(N720), .S(N719), .A(N476), .B(N452), .CI(N426));
ADDFX1 inst_cellmath__198_0_I322 (.CO(N722), .S(N721), .A(N454), .B(N500), .CI(N478));
ADDFX1 inst_cellmath__198_0_I323 (.CO(N724), .S(N723), .A(N607), .B(N540), .CI(N502));
ADDHX1 inst_cellmath__198_0_I324 (.CO(N726), .S(N725), .A(N110), .B(N230));
ADDHX1 inst_cellmath__198_0_I325 (.CO(N728), .S(N727), .A(N154), .B(N112));
ADDFX1 inst_cellmath__198_0_I326 (.CO(N730), .S(N729), .A(N270), .B(N156), .CI(N196));
ADDFX1 inst_cellmath__198_0_I327 (.CO(N732), .S(N731), .A(N198), .B(N116), .CI(N658));
ADDFX1 inst_cellmath__198_0_I328 (.CO(N734), .S(N733), .A(N660), .B(N200), .CI(N663));
ADDFX1 inst_cellmath__198_0_I329 (.CO(N736), .S(N735), .A(N662), .B(N664), .CI(N667));
ADDFX1 inst_cellmath__198_0_I330 (.CO(N738), .S(N737), .A(N666), .B(N668), .CI(N669));
ADDFX1 inst_cellmath__198_0_I331 (.CO(N740), .S(N739), .A(N673), .B(N670), .CI(N672));
ADDFX1 inst_cellmath__198_0_I332 (.CO(N742), .S(N741), .A(N676), .B(N674), .CI(N677));
ADDFX1 inst_cellmath__198_0_I333 (.CO(N744), .S(N743), .A(N681), .B(N678), .CI(N680));
ADDFX1 inst_cellmath__198_0_I334 (.CO(N746), .S(N745), .A(N684), .B(N682), .CI(N685));
ADDFX1 inst_cellmath__198_0_I335 (.CO(N748), .S(N747), .A(N689), .B(N686), .CI(N688));
ADDFX1 inst_cellmath__198_0_I336 (.CO(N750), .S(N749), .A(N693), .B(N690), .CI(N692));
ADDFX1 inst_cellmath__198_0_I337 (.CO(N752), .S(N751), .A(N697), .B(N694), .CI(N696));
ADDFX1 inst_cellmath__198_0_I338 (.CO(N754), .S(N753), .A(N701), .B(N698), .CI(N700));
ADDFX1 inst_cellmath__198_0_I339 (.CO(N756), .S(N755), .A(N705), .B(N702), .CI(N704));
ADDFX1 inst_cellmath__198_0_I340 (.CO(N758), .S(N757), .A(N709), .B(N706), .CI(N708));
ADDFX1 inst_cellmath__198_0_I341 (.CO(N760), .S(N759), .A(N713), .B(N710), .CI(N712));
ADDFX1 inst_cellmath__198_0_I342 (.CO(N762), .S(N761), .A(N717), .B(N714), .CI(N719));
ADDFX1 inst_cellmath__198_0_I343 (.CO(N764), .S(N763), .A(N718), .B(N606), .CI(N720));
ADDFX1 inst_cellmath__198_0_I344 (.CO(N766), .S(N765), .A(N480), .B(N522), .CI(N722));
ADDFX1 inst_cellmath__198_0_I345 (.CO(N768), .S(N767), .A(N524), .B(N504), .CI(N608));
ADDFX1 inst_cellmath__198_0_I346 (.CO(N770), .S(N769), .A(N609), .B(N560), .CI(N544));
ADDHX1 inst_cellmath__198_0_I347 (.CO(N772), .S(N771), .A(N106), .B(N148));
ADDHX1 inst_cellmath__198_0_I348 (.CO(N774), .S(N773), .A(N150), .B(N108));
ADDFX1 inst_cellmath__198_0_I349 (.CO(N776), .S(N775), .A(N192), .B(N152), .CI(N725));
ADDFX1 inst_cellmath__198_0_I350 (.CO(N778), .S(N777), .A(N726), .B(N194), .CI(N727));
ADDFX1 inst_cellmath__198_0_I351 (.CO(N780), .S(N779), .A(N657), .B(N728), .CI(N729));
ADDFX1 inst_cellmath__198_0_I352 (.CO(N782), .S(N781), .A(N730), .B(N659), .CI(N731));
ADDFX1 inst_cellmath__198_0_I353 (.CO(N784), .S(N783), .A(N661), .B(N732), .CI(N733));
ADDFX1 inst_cellmath__198_0_I354 (.CO(N786), .S(N785), .A(N734), .B(N665), .CI(N735));
ADDFX1 inst_cellmath__198_0_I355 (.CO(N788), .S(N787), .A(N671), .B(N736), .CI(N737));
ADDFX1 inst_cellmath__198_0_I356 (.CO(N790), .S(N789), .A(N738), .B(N675), .CI(N739));
ADDFX1 inst_cellmath__198_0_I357 (.CO(N792), .S(N791), .A(N679), .B(N740), .CI(N741));
ADDFX1 inst_cellmath__198_0_I358 (.CO(N794), .S(N793), .A(N683), .B(N742), .CI(N743));
ADDFX1 inst_cellmath__198_0_I359 (.CO(N796), .S(N795), .A(N744), .B(N687), .CI(N745));
ADDFX1 inst_cellmath__198_0_I360 (.CO(N798), .S(N797), .A(N746), .B(N691), .CI(N747));
ADDFX1 inst_cellmath__198_0_I361 (.CO(N800), .S(N799), .A(N748), .B(N695), .CI(N749));
ADDFX1 inst_cellmath__198_0_I362 (.CO(N802), .S(N801), .A(N750), .B(N699), .CI(N751));
ADDFX1 inst_cellmath__198_0_I363 (.CO(N804), .S(N803), .A(N752), .B(N703), .CI(N753));
ADDFX1 inst_cellmath__198_0_I364 (.CO(N806), .S(N805), .A(N754), .B(N707), .CI(N755));
ADDFX1 inst_cellmath__198_0_I365 (.CO(N808), .S(N807), .A(N756), .B(N711), .CI(N757));
ADDFX1 inst_cellmath__198_0_I366 (.CO(N810), .S(N809), .A(N758), .B(N715), .CI(N759));
ADDFX1 inst_cellmath__198_0_I367 (.CO(N812), .S(N811), .A(N761), .B(N716), .CI(N760));
ADDFX1 inst_cellmath__198_0_I368 (.CO(N814), .S(N813), .A(N763), .B(N721), .CI(N762));
ADDFX1 inst_cellmath__198_0_I369 (.CO(N816), .S(N815), .A(N764), .B(N723), .CI(N765));
ADDFX1 inst_cellmath__198_0_I370 (.CO(N818), .S(N817), .A(N767), .B(N724), .CI(N766));
ADDFX1 inst_cellmath__198_0_I371 (.CO(N820), .S(N819), .A(N768), .B(N526), .CI(N769));
ADDFX1 inst_cellmath__198_0_I372 (.CO(N822), .S(N821), .A(N610), .B(N546), .CI(N770));
ADDFX1 inst_cellmath__198_0_I373 (.CO(N824), .S(N823), .A(N611), .B(N578), .CI(N564));
NOR2XL inst_cellmath__198_0_I374 (.Y(N825), .A(N102), .B(N1577));
NOR2XL inst_cellmath__198_0_I376 (.Y(N827), .A(N188), .B(N771));
NAND2XL inst_cellmath__198_0_I377 (.Y(N828), .A(N188), .B(N771));
NOR2XL inst_cellmath__198_0_I378 (.Y(N829), .A(N772), .B(N773));
NAND2XL inst_cellmath__198_0_I379 (.Y(N830), .A(N772), .B(N773));
NOR2XL inst_cellmath__198_0_I380 (.Y(N831), .A(N774), .B(N775));
NAND2XL inst_cellmath__198_0_I381 (.Y(N832), .A(N774), .B(N775));
NOR2XL inst_cellmath__198_0_I382 (.Y(N833), .A(N776), .B(N777));
NAND2XL inst_cellmath__198_0_I383 (.Y(N834), .A(N776), .B(N777));
NOR2XL inst_cellmath__198_0_I384 (.Y(N835), .A(N778), .B(N779));
NAND2XL inst_cellmath__198_0_I385 (.Y(N836), .A(N778), .B(N779));
NOR2XL inst_cellmath__198_0_I386 (.Y(N837), .A(N780), .B(N781));
NAND2XL inst_cellmath__198_0_I387 (.Y(N838), .A(N780), .B(N781));
NOR2XL inst_cellmath__198_0_I388 (.Y(N839), .A(N782), .B(N783));
NAND2XL inst_cellmath__198_0_I389 (.Y(N840), .A(N782), .B(N783));
NOR2XL inst_cellmath__198_0_I390 (.Y(N841), .A(N784), .B(N785));
NAND2XL inst_cellmath__198_0_I391 (.Y(N842), .A(N784), .B(N785));
AND2XL inst_cellmath__198_0_I394 (.Y(N845), .A(N826), .B(N825));
INVXL inst_cellmath__198_0_I969 (.Y(N1594), .A(N827));
INVXL inst_cellmath__198_0_I970 (.Y(N1595), .A(N828));
OAI21XL inst_cellmath__198_0_I402 (.Y(N855), .A0(N1595), .A1(N845), .B0(N1594));
AOI21XL inst_cellmath__198_0_I410 (.Y(N863), .A0(N830), .A1(N855), .B0(N829));
INVXL inst_cellmath__198_0_I976 (.Y(N1601), .A(N831));
INVXL inst_cellmath__198_0_I977 (.Y(N1602), .A(N832));
OAI21XL inst_cellmath__198_0_I422 (.Y(N875), .A0(N1602), .A1(N863), .B0(N1601));
AOI21XL inst_cellmath__198_0_I434 (.Y(N887), .A0(N834), .A1(N875), .B0(N833));
INVXL inst_cellmath__198_0_I987 (.Y(N1612), .A(N835));
INVXL inst_cellmath__198_0_I988 (.Y(N1613), .A(N836));
OAI21XL inst_cellmath__198_0_I450 (.Y(N903), .A0(N1613), .A1(N887), .B0(N1612));
AOI21XL inst_cellmath__198_0_I466 (.Y(N919), .A0(N838), .A1(N903), .B0(N837));
INVXL inst_cellmath__198_0_I1004 (.Y(N1629), .A(N839));
INVXL inst_cellmath__198_0_I1005 (.Y(N1630), .A(N840));
AOI21XL inst_cellmath__198_0_I470 (.Y(N923), .A0(N842), .A1(N839), .B0(N841));
NAND2XL inst_cellmath__198_0_I471 (.Y(N924), .A(N842), .B(N840));
OAI21XL inst_cellmath__198_0_I488 (.Y(N941), .A0(N1630), .A1(N919), .B0(N1629));
OAI21XL inst_cellmath__198_0_I490 (.Y(N988), .A0(N924), .A1(N919), .B0(N923));
NAND2BXL inst_cellmath__198_0_I500 (.Y(N955), .AN(N827), .B(N828));
NAND2BXL inst_cellmath__198_0_I503 (.Y(N958), .AN(N829), .B(N830));
NAND2BXL inst_cellmath__198_0_I506 (.Y(N961), .AN(N831), .B(N832));
NAND2BXL inst_cellmath__198_0_I509 (.Y(N964), .AN(N833), .B(N834));
NAND2BXL inst_cellmath__198_0_I512 (.Y(N967), .AN(N835), .B(N836));
NAND2BXL inst_cellmath__198_0_I515 (.Y(N970), .AN(N837), .B(N838));
NAND2BXL inst_cellmath__198_0_I518 (.Y(N973), .AN(N839), .B(N840));
NAND2BXL inst_cellmath__198_0_I521 (.Y(N976), .AN(N841), .B(N842));
XOR2XL inst_cellmath__198_0_I2152 (.Y(inst_cellmath__198_0_out0[2]), .A(N102), .B(N1577));
XOR2XL inst_cellmath__198_0_I1073 (.Y(inst_cellmath__198_0_out0[3]), .A(N825), .B(N826));
XNOR2X1 inst_cellmath__198_0_I944 (.Y(inst_cellmath__198_0_out0[4]), .A(N845), .B(N955));
XOR2XL inst_cellmath__198_0_I1074 (.Y(inst_cellmath__198_0_out0[5]), .A(N855), .B(N958));
XNOR2X1 inst_cellmath__198_0_I1053 (.Y(inst_cellmath__198_0_out0[6]), .A(N863), .B(N961));
XOR2XL inst_cellmath__198_0_I1054 (.Y(inst_cellmath__198_0_out0[7]), .A(N875), .B(N964));
XNOR2X1 inst_cellmath__198_0_I528 (.Y(inst_cellmath__198_0_out0[8]), .A(N887), .B(N967));
XOR2XL inst_cellmath__198_0_I1055 (.Y(inst_cellmath__198_0_out0[9]), .A(N903), .B(N970));
XNOR2X1 inst_cellmath__198_0_I530 (.Y(inst_cellmath__198_0_out0[10]), .A(N919), .B(N973));
XOR2XL inst_cellmath__198_0_I531 (.Y(inst_cellmath__198_0_out0[11]), .A(N941), .B(N976));
NOR2XL inst_cellmath__198_0_I534 (.Y(N990), .A(N786), .B(N787));
NAND2XL inst_cellmath__198_0_I535 (.Y(N991), .A(N786), .B(N787));
NOR2XL inst_cellmath__198_0_I536 (.Y(N992), .A(N788), .B(N789));
NAND2XL inst_cellmath__198_0_I537 (.Y(N993), .A(N788), .B(N789));
NOR2XL inst_cellmath__198_0_I538 (.Y(N994), .A(N790), .B(N791));
NAND2XL inst_cellmath__198_0_I539 (.Y(N995), .A(N790), .B(N791));
NOR2XL inst_cellmath__198_0_I540 (.Y(N996), .A(N792), .B(N793));
NAND2XL inst_cellmath__198_0_I541 (.Y(N997), .A(N792), .B(N793));
NOR2XL inst_cellmath__198_0_I542 (.Y(N998), .A(N794), .B(N795));
NAND2XL inst_cellmath__198_0_I543 (.Y(N999), .A(N794), .B(N795));
NOR2XL inst_cellmath__198_0_I544 (.Y(N1000), .A(N796), .B(N797));
NAND2XL inst_cellmath__198_0_I545 (.Y(N1001), .A(N796), .B(N797));
NOR2XL inst_cellmath__198_0_I546 (.Y(N1002), .A(N798), .B(N799));
NAND2XL inst_cellmath__198_0_I547 (.Y(N1003), .A(N798), .B(N799));
NOR2XL inst_cellmath__198_0_I548 (.Y(N1004), .A(N800), .B(N801));
NAND2XL inst_cellmath__198_0_I549 (.Y(N1005), .A(N800), .B(N801));
NOR2XL inst_cellmath__198_0_I550 (.Y(N1006), .A(N802), .B(N803));
NAND2XL inst_cellmath__198_0_I551 (.Y(N1007), .A(N802), .B(N803));
NOR2XL inst_cellmath__198_0_I552 (.Y(N1008), .A(N804), .B(N805));
NAND2XL inst_cellmath__198_0_I553 (.Y(N1009), .A(N804), .B(N805));
NOR2XL inst_cellmath__198_0_I554 (.Y(N1010), .A(N806), .B(N807));
NAND2XL inst_cellmath__198_0_I555 (.Y(N1011), .A(N806), .B(N807));
NOR2XL inst_cellmath__198_0_I556 (.Y(N1012), .A(N808), .B(N809));
NAND2XL inst_cellmath__198_0_I557 (.Y(N1013), .A(N808), .B(N809));
NOR2XL inst_cellmath__198_0_I558 (.Y(N1014), .A(N811), .B(N810));
NAND2XL inst_cellmath__198_0_I559 (.Y(N1015), .A(N811), .B(N810));
NOR2XL inst_cellmath__198_0_I560 (.Y(N1016), .A(N813), .B(N812));
NAND2XL inst_cellmath__198_0_I561 (.Y(N1017), .A(N813), .B(N812));
NOR2XL inst_cellmath__198_0_I562 (.Y(N1018), .A(N814), .B(N815));
NAND2XL inst_cellmath__198_0_I563 (.Y(N1019), .A(N814), .B(N815));
NOR2XL inst_cellmath__198_0_I564 (.Y(N1020), .A(N817), .B(N816));
NAND2XL inst_cellmath__198_0_I565 (.Y(N1021), .A(N817), .B(N816));
NOR2XL inst_cellmath__198_0_I566 (.Y(N1022), .A(N818), .B(N819));
NAND2XL inst_cellmath__198_0_I567 (.Y(N1023), .A(N818), .B(N819));
NOR2XL inst_cellmath__198_0_I568 (.Y(N1024), .A(N821), .B(N820));
NAND2XL inst_cellmath__198_0_I569 (.Y(N1025), .A(N821), .B(N820));
NOR2XL inst_cellmath__198_0_I570 (.Y(N1026), .A(N823), .B(N822));
NAND2XL inst_cellmath__198_0_I571 (.Y(N1027), .A(N823), .B(N822));
NOR2XL inst_cellmath__198_0_I572 (.Y(N1028), .A(N612), .B(N824));
NAND2XL inst_cellmath__198_0_I573 (.Y(N1029), .A(N612), .B(N824));
AO21XL inst_cellmath__198_0_I578 (.Y(N1034), .A0(N991), .A1(N988), .B0(N990));
AO21XL inst_cellmath__198_0_I580 (.Y(N1036), .A0(N993), .A1(N990), .B0(N992));
AND2XL inst_cellmath__198_0_I581 (.Y(N1037), .A(N993), .B(N991));
AO21XL inst_cellmath__198_0_I582 (.Y(N1038), .A0(N995), .A1(N992), .B0(N994));
AND2XL inst_cellmath__198_0_I583 (.Y(N1039), .A(N995), .B(N993));
AO21XL inst_cellmath__198_0_I584 (.Y(N1040), .A0(N997), .A1(N994), .B0(N996));
AND2XL inst_cellmath__198_0_I585 (.Y(N1041), .A(N997), .B(N995));
AO21XL inst_cellmath__198_0_I586 (.Y(N1042), .A0(N999), .A1(N996), .B0(N998));
AND2XL inst_cellmath__198_0_I587 (.Y(N1043), .A(N999), .B(N997));
AO21XL inst_cellmath__198_0_I588 (.Y(N1044), .A0(N1001), .A1(N998), .B0(N1000));
AND2XL inst_cellmath__198_0_I589 (.Y(N1045), .A(N1001), .B(N999));
AO21XL inst_cellmath__198_0_I590 (.Y(N1046), .A0(N1003), .A1(N1000), .B0(N1002));
AND2XL inst_cellmath__198_0_I591 (.Y(N1047), .A(N1003), .B(N1001));
AO21XL inst_cellmath__198_0_I592 (.Y(N1048), .A0(N1005), .A1(N1002), .B0(N1004));
AND2XL inst_cellmath__198_0_I593 (.Y(N1049), .A(N1005), .B(N1003));
AO21XL inst_cellmath__198_0_I594 (.Y(N1050), .A0(N1007), .A1(N1004), .B0(N1006));
AND2XL inst_cellmath__198_0_I595 (.Y(N1051), .A(N1007), .B(N1005));
AO21XL inst_cellmath__198_0_I596 (.Y(N1052), .A0(N1009), .A1(N1006), .B0(N1008));
AND2XL inst_cellmath__198_0_I597 (.Y(N1053), .A(N1009), .B(N1007));
AO21XL inst_cellmath__198_0_I598 (.Y(N1054), .A0(N1011), .A1(N1008), .B0(N1010));
AND2XL inst_cellmath__198_0_I599 (.Y(N1055), .A(N1011), .B(N1009));
AO21XL inst_cellmath__198_0_I600 (.Y(N1056), .A0(N1013), .A1(N1010), .B0(N1012));
AND2XL inst_cellmath__198_0_I601 (.Y(N1057), .A(N1013), .B(N1011));
AO21XL inst_cellmath__198_0_I602 (.Y(N1058), .A0(N1015), .A1(N1012), .B0(N1014));
AND2XL inst_cellmath__198_0_I603 (.Y(N1059), .A(N1015), .B(N1013));
AO21XL inst_cellmath__198_0_I604 (.Y(N1060), .A0(N1017), .A1(N1014), .B0(N1016));
AND2XL inst_cellmath__198_0_I605 (.Y(N1061), .A(N1017), .B(N1015));
AO21XL inst_cellmath__198_0_I606 (.Y(N1062), .A0(N1019), .A1(N1016), .B0(N1018));
AND2XL inst_cellmath__198_0_I607 (.Y(N1063), .A(N1019), .B(N1017));
AO21XL inst_cellmath__198_0_I608 (.Y(N1064), .A0(N1021), .A1(N1018), .B0(N1020));
AND2XL inst_cellmath__198_0_I609 (.Y(N1065), .A(N1021), .B(N1019));
AO21XL inst_cellmath__198_0_I610 (.Y(N1066), .A0(N1023), .A1(N1020), .B0(N1022));
AND2XL inst_cellmath__198_0_I611 (.Y(N1067), .A(N1023), .B(N1021));
AO21XL inst_cellmath__198_0_I612 (.Y(N1068), .A0(N1025), .A1(N1022), .B0(N1024));
AND2XL inst_cellmath__198_0_I613 (.Y(N1069), .A(N1025), .B(N1023));
AO21XL inst_cellmath__198_0_I614 (.Y(N1070), .A0(N1027), .A1(N1024), .B0(N1026));
AND2XL inst_cellmath__198_0_I615 (.Y(N1071), .A(N1027), .B(N1025));
AO21XL inst_cellmath__198_0_I616 (.Y(N1072), .A0(N1029), .A1(N1026), .B0(N1028));
AND2XL inst_cellmath__198_0_I617 (.Y(N1073), .A(N1029), .B(N1027));
AO21XL inst_cellmath__198_0_I624 (.Y(N1080), .A0(N988), .A1(N1037), .B0(N1036));
AO21XL inst_cellmath__198_0_I626 (.Y(N1082), .A0(N1039), .A1(N1034), .B0(N1038));
AO21XL inst_cellmath__198_0_I628 (.Y(N1084), .A0(N1041), .A1(N1036), .B0(N1040));
AND2XL inst_cellmath__198_0_I629 (.Y(N1085), .A(N1041), .B(N1037));
AO21XL inst_cellmath__198_0_I630 (.Y(N1086), .A0(N1043), .A1(N1038), .B0(N1042));
AND2XL inst_cellmath__198_0_I631 (.Y(N1087), .A(N1043), .B(N1039));
AO21XL inst_cellmath__198_0_I632 (.Y(N1088), .A0(N1045), .A1(N1040), .B0(N1044));
AND2XL inst_cellmath__198_0_I633 (.Y(N1089), .A(N1045), .B(N1041));
AO21XL inst_cellmath__198_0_I634 (.Y(N1090), .A0(N1047), .A1(N1042), .B0(N1046));
AND2XL inst_cellmath__198_0_I635 (.Y(N1091), .A(N1047), .B(N1043));
AO21XL inst_cellmath__198_0_I636 (.Y(N1092), .A0(N1049), .A1(N1044), .B0(N1048));
AND2XL inst_cellmath__198_0_I637 (.Y(N1093), .A(N1049), .B(N1045));
AO21XL inst_cellmath__198_0_I638 (.Y(N1094), .A0(N1051), .A1(N1046), .B0(N1050));
AND2XL inst_cellmath__198_0_I639 (.Y(N1095), .A(N1051), .B(N1047));
AO21XL inst_cellmath__198_0_I640 (.Y(N1096), .A0(N1053), .A1(N1048), .B0(N1052));
AND2XL inst_cellmath__198_0_I641 (.Y(N1097), .A(N1053), .B(N1049));
AO21XL inst_cellmath__198_0_I642 (.Y(N1098), .A0(N1055), .A1(N1050), .B0(N1054));
AND2XL inst_cellmath__198_0_I643 (.Y(N1099), .A(N1055), .B(N1051));
AO21XL inst_cellmath__198_0_I644 (.Y(N1100), .A0(N1057), .A1(N1052), .B0(N1056));
AND2XL inst_cellmath__198_0_I645 (.Y(N1101), .A(N1057), .B(N1053));
AO21XL inst_cellmath__198_0_I646 (.Y(N1102), .A0(N1059), .A1(N1054), .B0(N1058));
AND2XL inst_cellmath__198_0_I647 (.Y(N1103), .A(N1059), .B(N1055));
AO21XL inst_cellmath__198_0_I648 (.Y(N1104), .A0(N1061), .A1(N1056), .B0(N1060));
AND2XL inst_cellmath__198_0_I649 (.Y(N1105), .A(N1061), .B(N1057));
AO21XL inst_cellmath__198_0_I650 (.Y(N1106), .A0(N1063), .A1(N1058), .B0(N1062));
AND2XL inst_cellmath__198_0_I651 (.Y(N1107), .A(N1063), .B(N1059));
AO21XL inst_cellmath__198_0_I652 (.Y(N1108), .A0(N1065), .A1(N1060), .B0(N1064));
AND2XL inst_cellmath__198_0_I653 (.Y(N1109), .A(N1065), .B(N1061));
AO21XL inst_cellmath__198_0_I654 (.Y(N1110), .A0(N1067), .A1(N1062), .B0(N1066));
AND2XL inst_cellmath__198_0_I655 (.Y(N1111), .A(N1067), .B(N1063));
AO21XL inst_cellmath__198_0_I656 (.Y(N1112), .A0(N1069), .A1(N1064), .B0(N1068));
AND2XL inst_cellmath__198_0_I657 (.Y(N1113), .A(N1069), .B(N1065));
AO21XL inst_cellmath__198_0_I658 (.Y(N1114), .A0(N1071), .A1(N1066), .B0(N1070));
AND2XL inst_cellmath__198_0_I659 (.Y(N1115), .A(N1071), .B(N1067));
AO21XL inst_cellmath__198_0_I660 (.Y(N1116), .A0(N1073), .A1(N1068), .B0(N1072));
AND2XL inst_cellmath__198_0_I661 (.Y(N1117), .A(N1073), .B(N1069));
AO21XL inst_cellmath__198_0_I672 (.Y(N1128), .A0(N1085), .A1(N988), .B0(N1084));
AO21XL inst_cellmath__198_0_I674 (.Y(N1130), .A0(N1087), .A1(N1034), .B0(N1086));
AO21XL inst_cellmath__198_0_I676 (.Y(N1132), .A0(N1089), .A1(N1080), .B0(N1088));
AO21XL inst_cellmath__198_0_I678 (.Y(N1134), .A0(N1091), .A1(N1082), .B0(N1090));
AO21XL inst_cellmath__198_0_I680 (.Y(N1136), .A0(N1093), .A1(N1084), .B0(N1092));
AND2XL inst_cellmath__198_0_I681 (.Y(N1137), .A(N1093), .B(N1085));
AO21XL inst_cellmath__198_0_I682 (.Y(N1138), .A0(N1095), .A1(N1086), .B0(N1094));
AND2XL inst_cellmath__198_0_I683 (.Y(N1139), .A(N1095), .B(N1087));
AO21XL inst_cellmath__198_0_I684 (.Y(N1140), .A0(N1097), .A1(N1088), .B0(N1096));
AND2XL inst_cellmath__198_0_I685 (.Y(N1141), .A(N1097), .B(N1089));
AO21XL inst_cellmath__198_0_I686 (.Y(N1142), .A0(N1099), .A1(N1090), .B0(N1098));
AND2XL inst_cellmath__198_0_I687 (.Y(N1143), .A(N1099), .B(N1091));
AO21XL inst_cellmath__198_0_I688 (.Y(N1144), .A0(N1101), .A1(N1092), .B0(N1100));
AND2XL inst_cellmath__198_0_I689 (.Y(N1145), .A(N1101), .B(N1093));
AO21XL inst_cellmath__198_0_I690 (.Y(N1146), .A0(N1103), .A1(N1094), .B0(N1102));
AO21XL inst_cellmath__198_0_I692 (.Y(N1148), .A0(N1105), .A1(N1096), .B0(N1104));
AO21XL inst_cellmath__198_0_I694 (.Y(N1150), .A0(N1107), .A1(N1098), .B0(N1106));
AO21XL inst_cellmath__198_0_I696 (.Y(N1152), .A0(N1109), .A1(N1100), .B0(N1108));
AND2XL inst_cellmath__198_0_I697 (.Y(N1153), .A(N1109), .B(N1101));
AO21XL inst_cellmath__198_0_I698 (.Y(N1154), .A0(N1111), .A1(N1102), .B0(N1110));
AND2XL inst_cellmath__198_0_I699 (.Y(N1155), .A(N1111), .B(N1103));
AO21XL inst_cellmath__198_0_I700 (.Y(N1156), .A0(N1113), .A1(N1104), .B0(N1112));
AND2XL inst_cellmath__198_0_I701 (.Y(N1157), .A(N1113), .B(N1105));
AO21XL inst_cellmath__198_0_I702 (.Y(N1158), .A0(N1115), .A1(N1106), .B0(N1114));
AND2XL inst_cellmath__198_0_I703 (.Y(N1159), .A(N1115), .B(N1107));
AO21XL inst_cellmath__198_0_I704 (.Y(N1160), .A0(N1117), .A1(N1108), .B0(N1116));
AND2XL inst_cellmath__198_0_I705 (.Y(N1161), .A(N1117), .B(N1109));
AO21XL inst_cellmath__198_0_I740 (.Y(N1196), .A0(N1153), .A1(N1136), .B0(N1152));
AND2XL inst_cellmath__198_0_I741 (.Y(N1197), .A(N1153), .B(N1137));
AO21XL inst_cellmath__198_0_I742 (.Y(N1198), .A0(N1155), .A1(N1138), .B0(N1154));
AND2XL inst_cellmath__198_0_I743 (.Y(N1199), .A(N1155), .B(N1139));
AO21XL inst_cellmath__198_0_I744 (.Y(N1200), .A0(N1157), .A1(N1140), .B0(N1156));
AND2XL inst_cellmath__198_0_I745 (.Y(N1201), .A(N1157), .B(N1141));
AO21XL inst_cellmath__198_0_I746 (.Y(N1202), .A0(N1159), .A1(N1142), .B0(N1158));
AND2XL inst_cellmath__198_0_I747 (.Y(N1203), .A(N1159), .B(N1143));
AO21XL inst_cellmath__198_0_I748 (.Y(N1204), .A0(N1161), .A1(N1144), .B0(N1160));
AND2XL inst_cellmath__198_0_I749 (.Y(N1205), .A(N1161), .B(N1145));
AOI21XL inst_cellmath__198_0_I1056 (.Y(N1668), .A0(N1137), .A1(N988), .B0(N1136));
AOI21XL inst_cellmath__198_0_I1057 (.Y(N1669), .A0(N1139), .A1(N1034), .B0(N1138));
AOI21XL inst_cellmath__198_0_I1058 (.Y(N1670), .A0(N1141), .A1(N1080), .B0(N1140));
AOI21XL inst_cellmath__198_0_I1059 (.Y(N1671), .A0(N1143), .A1(N1082), .B0(N1142));
AOI21XL inst_cellmath__198_0_I1060 (.Y(N1672), .A0(N1145), .A1(N1128), .B0(N1144));
AOI31X1 inst_cellmath__198_0_I1075 (.Y(N1673), .A0(N1103), .A1(N1095), .A2(N1130), .B0(N1146));
AOI31X1 inst_cellmath__198_0_I1076 (.Y(N1674), .A0(N1105), .A1(N1097), .A2(N1132), .B0(N1148));
AOI31X1 inst_cellmath__198_0_I1077 (.Y(N1675), .A0(N1107), .A1(N1099), .A2(N1134), .B0(N1150));
AO21XL inst_cellmath__198_0_I784 (.Y(N1240), .A0(N1197), .A1(N988), .B0(N1196));
AO21XL inst_cellmath__198_0_I786 (.Y(N1242), .A0(N1199), .A1(N1034), .B0(N1198));
AO21XL inst_cellmath__198_0_I788 (.Y(N1244), .A0(N1201), .A1(N1080), .B0(N1200));
AO21XL inst_cellmath__198_0_I790 (.Y(N1246), .A0(N1203), .A1(N1082), .B0(N1202));
AO21XL inst_cellmath__198_0_I792 (.Y(N1248), .A0(N1205), .A1(N1128), .B0(N1204));
NAND2BXL inst_cellmath__198_0_I801 (.Y(N1257), .AN(N990), .B(N991));
NAND2BXL inst_cellmath__198_0_I804 (.Y(N1260), .AN(N992), .B(N993));
NAND2BXL inst_cellmath__198_0_I807 (.Y(N1263), .AN(N994), .B(N995));
NAND2BXL inst_cellmath__198_0_I810 (.Y(N1266), .AN(N996), .B(N997));
NAND2BXL inst_cellmath__198_0_I813 (.Y(N1269), .AN(N998), .B(N999));
NAND2BXL inst_cellmath__198_0_I816 (.Y(N1272), .AN(N1000), .B(N1001));
NAND2BXL inst_cellmath__198_0_I819 (.Y(N1275), .AN(N1002), .B(N1003));
NAND2BXL inst_cellmath__198_0_I822 (.Y(N1278), .AN(N1004), .B(N1005));
NAND2BXL inst_cellmath__198_0_I825 (.Y(N1281), .AN(N1006), .B(N1007));
NAND2BXL inst_cellmath__198_0_I828 (.Y(N1284), .AN(N1008), .B(N1009));
NAND2BXL inst_cellmath__198_0_I831 (.Y(N1287), .AN(N1010), .B(N1011));
NAND2BXL inst_cellmath__198_0_I834 (.Y(N1290), .AN(N1012), .B(N1013));
NAND2BXL inst_cellmath__198_0_I837 (.Y(N1293), .AN(N1014), .B(N1015));
NAND2BXL inst_cellmath__198_0_I840 (.Y(N1296), .AN(N1016), .B(N1017));
NAND2BXL inst_cellmath__198_0_I843 (.Y(N1299), .AN(N1018), .B(N1019));
NAND2BXL inst_cellmath__198_0_I846 (.Y(N1302), .AN(N1020), .B(N1021));
NAND2BXL inst_cellmath__198_0_I849 (.Y(N1305), .AN(N1022), .B(N1023));
NAND2BXL inst_cellmath__198_0_I852 (.Y(N1308), .AN(N1024), .B(N1025));
NAND2BXL inst_cellmath__198_0_I855 (.Y(N1311), .AN(N1026), .B(N1027));
NAND2BXL inst_cellmath__198_0_I858 (.Y(N1314), .AN(N1028), .B(N1029));
NOR2BX1 inst_cellmath__198_0_I1079 (.Y(N1317), .AN(N1591), .B(N1592));
XOR2XL inst_cellmath__198_0_I1065 (.Y(inst_cellmath__198_0_out0[12]), .A(N988), .B(N1257));
XOR2XL inst_cellmath__198_0_I1066 (.Y(inst_cellmath__198_0_out0[13]), .A(N1034), .B(N1260));
XOR2XL inst_cellmath__198_0_I1067 (.Y(inst_cellmath__198_0_out0[14]), .A(N1080), .B(N1263));
XOR2XL inst_cellmath__198_0_I1068 (.Y(inst_cellmath__198_0_out0[15]), .A(N1082), .B(N1266));
XOR2XL inst_cellmath__198_0_I1069 (.Y(inst_cellmath__198_0_out0[16]), .A(N1128), .B(N1269));
XOR2XL inst_cellmath__198_0_I1070 (.Y(inst_cellmath__198_0_out0[17]), .A(N1130), .B(N1272));
XOR2XL inst_cellmath__198_0_I1071 (.Y(inst_cellmath__198_0_out0[18]), .A(N1132), .B(N1275));
XOR2XL inst_cellmath__198_0_I1072 (.Y(inst_cellmath__198_0_out0[19]), .A(N1134), .B(N1278));
XNOR2X1 inst_cellmath__198_0_I871 (.Y(inst_cellmath__198_0_out0[20]), .A(N1668), .B(N1281));
XNOR2X1 inst_cellmath__198_0_I872 (.Y(inst_cellmath__198_0_out0[21]), .A(N1669), .B(N1284));
XNOR2X1 inst_cellmath__198_0_I873 (.Y(inst_cellmath__198_0_out0[22]), .A(N1670), .B(N1287));
XNOR2X1 inst_cellmath__198_0_I874 (.Y(inst_cellmath__198_0_out0[23]), .A(N1671), .B(N1290));
XNOR2X1 inst_cellmath__198_0_I875 (.Y(inst_cellmath__198_0_out0[24]), .A(N1672), .B(N1293));
XNOR2X1 inst_cellmath__198_0_I876 (.Y(inst_cellmath__198_0_out0[25]), .A(N1673), .B(N1296));
XNOR2X1 inst_cellmath__198_0_I877 (.Y(inst_cellmath__198_0_out0[26]), .A(N1674), .B(N1299));
XNOR2X1 inst_cellmath__198_0_I878 (.Y(inst_cellmath__198_0_out0[27]), .A(N1675), .B(N1302));
XOR2XL inst_cellmath__198_0_I879 (.Y(inst_cellmath__198_0_out0[28]), .A(N1240), .B(N1305));
XOR2XL inst_cellmath__198_0_I880 (.Y(inst_cellmath__198_0_out0[29]), .A(N1242), .B(N1308));
XOR2XL inst_cellmath__198_0_I881 (.Y(inst_cellmath__198_0_out0[30]), .A(N1244), .B(N1311));
XOR2XL inst_cellmath__198_0_I882 (.Y(inst_cellmath__198_0_out0[31]), .A(N1246), .B(N1314));
XOR2XL inst_cellmath__198_0_I883 (.Y(inst_cellmath__198_0_out0[32]), .A(N1248), .B(N1317));
assign inst_cellmath__198_0_out0[1] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__203_0_bdw1114505291_bdw (
	inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1,
	inst_cellmath__203_0_in0,
	inst_cellmath__203_0_in1,
	inst_cellmath__203_0_in2,
	inst_cellmath__203_0_in3,
	inst_cellmath__203_0_in4
	); /* architecture "gate_level" */ 
output [46:0] inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1;
input [15:0] inst_cellmath__203_0_in0;
input [32:17] inst_cellmath__203_0_in1;
input [42:23] inst_cellmath__203_0_in2;
input [21:0] inst_cellmath__203_0_in3;
input [0:0] inst_cellmath__203_0_in4;
wire N518,N520,N522,N524,N526,N528,N530 
	,N532,N534,N536,N538,N540,N542,N544,N546 
	,N548,N550,N552,N554,N566,N567,N568,N569 
	,N570,N571,N572,N573,N574,N575,N576,N577 
	,N578,N579,N580,N581,N582,N583,N584,N585 
	,N588,N589,N595,N596,N597,N598,N599,N600 
	,N601,N602,N603,N604,N605,N606,N607,N608 
	,N609,N610,N611,N612,N613,N614,N615,N618 
	,N619,N625,N626,N627,N628,N629,N630,N631 
	,N632,N633,N634,N635,N636,N637,N638,N639 
	,N640,N641,N642,N643,N644,N645,N648,N649 
	,N655,N656,N657,N658,N659,N660,N661,N662 
	,N663,N664,N665,N666,N667,N668,N669,N670 
	,N671,N672,N673,N674,N675,N678,N679,N685 
	,N686,N687,N688,N689,N690,N691,N692,N693 
	,N694,N695,N696,N697,N698,N699,N700,N701 
	,N702,N703,N704,N705,N708,N709,N715,N716 
	,N717,N718,N719,N720,N721,N722,N723,N724 
	,N725,N726,N727,N728,N729,N730,N731,N732 
	,N733,N734,N735,N738,N739,N745,N746,N747 
	,N748,N749,N750,N751,N752,N753,N754,N755 
	,N756,N757,N758,N759,N760,N761,N762,N763 
	,N764,N765,N768,N770,N779,N781,N783,N785 
	,N787,N789,N791,N793,N795,N797,N799,N801 
	,N803,N805,N807,N809,N811,N813,N815,N817 
	,N819,N1025,N1027,N1029,N1031,N1033,N1035,N1037 
	,N1039,N1041,N1043,N1045,N1047,N1049,N1051,N1053 
	,N1055,N1059,N1061,N1067,N1077,N1078,N1079,N1080 
	,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088 
	,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096 
	,N1097,N1098,N1099,N1102,N1103,N1109,N1110,N1111 
	,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119 
	,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127 
	,N1128,N1129,N1130,N1131,N1134,N1135,N1141,N1142 
	,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150 
	,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158 
	,N1159,N1160,N1161,N1162,N1163,N1166,N1167,N1173 
	,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181 
	,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189 
	,N1190,N1191,N1192,N1193,N1194,N1195,N1198,N1199 
	,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212 
	,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220 
	,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1230 
	,N1231,N1237,N1238,N1239,N1240,N1241,N1242,N1243 
	,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251 
	,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259 
	,N1262,N1263,N1269,N1270,N1271,N1272,N1273,N1274 
	,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282 
	,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290 
	,N1294,N1295,N1301,N1302,N1303,N1304,N1305,N1306 
	,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314 
	,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322 
	,N1366,N1379,N1380,N1383,N1384,N1387,N1388,N1389 
	,N1390,N1391,N1392,N1395,N1396,N1397,N1398,N1399 
	,N1400,N1403,N1404,N1405,N1406,N1407,N1408,N1409 
	,N1410,N1411,N1412,N1415,N1416,N1417,N1418,N1419 
	,N1420,N1421,N1422,N1423,N1424,N1427,N1428,N1429 
	,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437 
	,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447 
	,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455 
	,N1456,N1459,N1460,N1461,N1462,N1463,N1464,N1465 
	,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473 
	,N1474,N1475,N1476,N1479,N1480,N1481,N1482,N1483 
	,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491 
	,N1492,N1493,N1494,N1495,N1496,N1499,N1500,N1501 
	,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509 
	,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517 
	,N1518,N1519,N1520,N1523,N1524,N1525,N1526,N1527 
	,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535 
	,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543 
	,N1544,N1547,N1548,N1549,N1550,N1551,N1552,N1553 
	,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561 
	,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569 
	,N1570,N1571,N1572,N1575,N1576,N1577,N1578,N1579 
	,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587 
	,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595 
	,N1596,N1597,N1598,N1599,N1600,N1603,N1604,N1605 
	,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613 
	,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621 
	,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629 
	,N1630,N1633,N1634,N1635,N1636,N1637,N1638,N1639 
	,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647 
	,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655 
	,N1656,N1657,N1658,N1659,N1660,N1663,N1664,N1665 
	,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673 
	,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681 
	,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689 
	,N1690,N1691,N1692,N1695,N1696,N1699,N1700,N1701 
	,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709 
	,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717 
	,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725 
	,N1726,N1729,N1730,N1732,N1733,N1734,N1735,N1736 
	,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744 
	,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752 
	,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760 
	,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770 
	,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778 
	,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786 
	,N1787,N1788,N1789,N1790,N1791,N1792,N1795,N1796 
	,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805 
	,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813 
	,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821 
	,N1822,N1823,N1824,N1827,N1828,N1830,N1831,N1832 
	,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840 
	,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848 
	,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856 
	,N1859,N1860,N1863,N1864,N1865,N1866,N1867,N1868 
	,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876 
	,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884 
	,N1885,N1886,N1887,N1888,N1891,N1892,N1893,N1894 
	,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902 
	,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910 
	,N1911,N1912,N1913,N1914,N1915,N1916,N1919,N1920 
	,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930 
	,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938 
	,N1939,N1940,N1941,N1942,N1943,N1944,N1947,N1948 
	,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958 
	,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966 
	,N1967,N1968,N1969,N1970,N1973,N1974,N1975,N1976 
	,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984 
	,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992 
	,N1995,N1996,N1999,N2000,N2001,N2002,N2003,N2004 
	,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012 
	,N2013,N2014,N2017,N2018,N2019,N2020,N2021,N2022 
	,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030 
	,N2031,N2032,N2035,N2036,N2039,N2040,N2041,N2042 
	,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050 
	,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060 
	,N2061,N2062,N2063,N2064,N2067,N2068,N2071,N2072 
	,N2073,N2074,N2075,N2076,N2077,N2078,N2081,N2082 
	,N2083,N2084,N2085,N2086,N2087,N2088,N2091,N2092 
	,N2095,N2096,N2097,N2098,N2101,N2102,N2103,N2104 
	,N2107,N2108,N2111,N2112,N2300,N2309,N2318,N2327 
	,N2336,N2345,N2354,N2363,N2372,N2381,N2390,N2399 
	,N2408,N2417,N2426,N2435,N2444,N2453,N2462,N2471 
	,N2480,N2491,N2502,N2511,N2520,N2529,N2538,N2547 
	,N2556,N2565,N2574,N2583,N2592,N2601,N2610,N2619 
	,N2628,N2637,N2646,N2655,N2664,N2673,N2682,N2693 
	,N2704,N2713,N2722,N2731,N2740,N2749,N2758,N2767 
	,N2776,N2785,N2794,N2803,N2812,N2821,N2830,N2839 
	,N2848,N2857,N2866,N2875,N2884,N2895,N2906,N2915 
	,N2924,N2933,N2942,N2951,N2960,N2969,N2978,N2987 
	,N2996,N3005,N3014,N3023,N3032,N3041,N3050,N3059 
	,N3068,N3077,N3086,N3097,N3108,N3117,N3126,N3135 
	,N3144,N3153,N3162,N3171,N3180,N3189,N3198,N3207 
	,N3216,N3225,N3234,N3243,N3252,N3261,N3270,N3279 
	,N3288,N3299,N3310,N3319,N3328,N3337,N3346,N3355 
	,N3364,N3373,N3382,N3391,N3400,N3409,N3418,N3427 
	,N3436,N3445,N3454,N3463,N3472,N3481,N3490,N3501 
	,N3512,N3521,N3530,N3539,N3548,N3557,N3566,N3575 
	,N3584,N3593,N3602,N3611,N3620,N3629,N3638,N3647 
	,N3656,N3665,N3674,N3683,N3692,N3714,N3723,N3732 
	,N3741,N3750,N3759,N3768,N3777,N3786,N3795,N3804 
	,N3813,N3822,N3831,N3840,N3849,N3858,N3867,N3876 
	,N3885,N3894,N3903,N3912,N3923,N3934,N3943,N3952 
	,N3961,N3970,N3979,N3988,N3997,N4006,N4015,N4024 
	,N4033,N4042,N4051,N4060,N4069,N4078,N4087,N4096 
	,N4105,N4114,N4123,N4132,N4143,N4154,N4163,N4172 
	,N4181,N4190,N4199,N4208,N4217,N4226,N4235,N4244 
	,N4253,N4262,N4271,N4280,N4289,N4298,N4307,N4316 
	,N4325,N4334,N4343,N4352,N4363,N4374,N4383,N4392 
	,N4401,N4410,N4419,N4428,N4437,N4446,N4455,N4464 
	,N4473,N4482,N4491,N4500,N4509,N4518,N4527,N4536 
	,N4545,N4554,N4563,N4572,N4583,N4594,N4603,N4612 
	,N4621,N4630,N4639,N4648,N4657,N4666,N4675,N4684 
	,N4693,N4702,N4711,N4720,N4729,N4738,N4747,N4756 
	,N4765,N4774,N4783,N4792,N4803,N4814,N4823,N4832 
	,N4841,N4850,N4859,N4868,N4877,N4886,N4895,N4904 
	,N4913,N4922,N4931,N4940,N4949,N4958,N4967,N4976 
	,N4985,N4994,N5003,N5012,N5023,N5034,N5043,N5052 
	,N5061,N5070,N5079,N5088,N5097,N5106,N5115,N5124 
	,N5133,N5142,N5151,N5160,N5169,N5178,N5187,N5196 
	,N5205,N5214,N5223,N5232,N5243,N5254,N5263,N5272 
	,N5281,N5290,N5299,N5308,N5317,N5326,N5335,N5344 
	,N5353,N5362,N5371,N5380,N5389,N5398,N5407,N5416 
	,N5425,N5434,N5443,N5452,N5461,N5479,N5488,N5509 
	,N5518,N5527,N5536,N5545,N5635,N5636,N5637,N5638 
	,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646 
	,N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654 
	,N5655,N5658,N5659,N5660,N5661,N5664,N5665,N5666 
	,N5669,N5670,N5671,N5674,N5675,N5676,N5679,N5680 
	,N5681,N5684,N5685,N5686,N5689,N5690,N5691,N5692 
	,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700 
	,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708 
	,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5718 
	,N5719,N5720,N5721,N5724,N5725,N5726,N5729,N5730 
	,N5731,N5734,N5735,N5736,N5739,N5740,N5741,N5744 
	,N5745,N5746,N5749,N5750,N5751,N5754;
INVXL inst_cellmath__203_0_I1839 (.Y(N5635), .A(inst_cellmath__203_0_in2[23]));
INVXL inst_cellmath__203_0_I1840 (.Y(N5636), .A(inst_cellmath__203_0_in2[24]));
INVXL inst_cellmath__203_0_I1841 (.Y(N5637), .A(inst_cellmath__203_0_in2[25]));
INVXL inst_cellmath__203_0_I1842 (.Y(N5638), .A(inst_cellmath__203_0_in2[26]));
INVXL inst_cellmath__203_0_I1843 (.Y(N5639), .A(inst_cellmath__203_0_in2[27]));
INVXL inst_cellmath__203_0_I1844 (.Y(N5640), .A(inst_cellmath__203_0_in2[28]));
INVXL inst_cellmath__203_0_I1845 (.Y(N5641), .A(inst_cellmath__203_0_in2[29]));
INVXL inst_cellmath__203_0_I1846 (.Y(N5642), .A(inst_cellmath__203_0_in2[30]));
INVXL inst_cellmath__203_0_I1847 (.Y(N5643), .A(inst_cellmath__203_0_in2[31]));
INVXL inst_cellmath__203_0_I1848 (.Y(N5644), .A(inst_cellmath__203_0_in2[32]));
INVXL inst_cellmath__203_0_I1849 (.Y(N5645), .A(inst_cellmath__203_0_in2[33]));
INVXL inst_cellmath__203_0_I1850 (.Y(N5646), .A(inst_cellmath__203_0_in2[34]));
INVXL inst_cellmath__203_0_I1851 (.Y(N5647), .A(inst_cellmath__203_0_in2[35]));
INVXL inst_cellmath__203_0_I1852 (.Y(N5648), .A(inst_cellmath__203_0_in2[36]));
INVXL inst_cellmath__203_0_I1853 (.Y(N5649), .A(inst_cellmath__203_0_in2[37]));
INVXL inst_cellmath__203_0_I1854 (.Y(N5650), .A(inst_cellmath__203_0_in2[38]));
INVXL inst_cellmath__203_0_I1855 (.Y(N5651), .A(inst_cellmath__203_0_in2[39]));
INVXL inst_cellmath__203_0_I1856 (.Y(N5652), .A(inst_cellmath__203_0_in2[40]));
INVXL inst_cellmath__203_0_I1857 (.Y(N5653), .A(inst_cellmath__203_0_in2[41]));
INVXL inst_cellmath__203_0_I1858 (.Y(N5654), .A(inst_cellmath__203_0_in2[42]));
INVXL inst_cellmath__203_0_I1859 (.Y(N5655), .A(inst_cellmath__203_0_in1[17]));
NOR2XL inst_cellmath__203_0_I71 (.Y(inst_cellmath__203_0_out1[0]), .A(N5655), .B(N5635));
NOR2XL inst_cellmath__203_0_I72 (.Y(N518), .A(N5655), .B(N5636));
NOR2XL inst_cellmath__203_0_I73 (.Y(N520), .A(N5655), .B(N5637));
NOR2XL inst_cellmath__203_0_I74 (.Y(N522), .A(N5655), .B(N5638));
NOR2XL inst_cellmath__203_0_I75 (.Y(N524), .A(N5655), .B(N5639));
NOR2XL inst_cellmath__203_0_I76 (.Y(N526), .A(N5655), .B(N5640));
NOR2XL inst_cellmath__203_0_I77 (.Y(N528), .A(N5655), .B(N5641));
NOR2XL inst_cellmath__203_0_I78 (.Y(N530), .A(N5655), .B(N5642));
NOR2XL inst_cellmath__203_0_I79 (.Y(N532), .A(N5655), .B(N5643));
NOR2XL inst_cellmath__203_0_I80 (.Y(N534), .A(N5655), .B(N5644));
NOR2XL inst_cellmath__203_0_I81 (.Y(N536), .A(N5655), .B(N5645));
NOR2XL inst_cellmath__203_0_I82 (.Y(N538), .A(N5655), .B(N5646));
NOR2XL inst_cellmath__203_0_I83 (.Y(N540), .A(N5655), .B(N5647));
NOR2XL inst_cellmath__203_0_I84 (.Y(N542), .A(N5655), .B(N5648));
NOR2XL inst_cellmath__203_0_I85 (.Y(N544), .A(N5655), .B(N5649));
NOR2XL inst_cellmath__203_0_I86 (.Y(N546), .A(N5655), .B(N5650));
NOR2XL inst_cellmath__203_0_I87 (.Y(N548), .A(N5655), .B(N5651));
NOR2XL inst_cellmath__203_0_I88 (.Y(N550), .A(N5655), .B(N5652));
NOR2XL inst_cellmath__203_0_I89 (.Y(N552), .A(N5655), .B(N5653));
NOR2XL inst_cellmath__203_0_I90 (.Y(N554), .A(N5655), .B(N5654));
INVXL inst_cellmath__203_0_I1862 (.Y(N5658), .A(inst_cellmath__203_0_in1[18]));
NAND2BX1 inst_cellmath__203_0_I1968 (.Y(N5659), .AN(inst_cellmath__203_0_in1[19]), .B(inst_cellmath__203_0_in1[18]));
INVXL inst_cellmath__203_0_I1864 (.Y(N5660), .A(inst_cellmath__203_0_in1[19]));
NOR2XL addgen2_A_I1066 (.Y(N2300), .A(N5635), .B(N5658));
MXI2XL addgen2_A_I1067 (.Y(inst_cellmath__203_0_out1[1]), .A(N5660), .B(N5659), .S0(N2300));
MXI2XL addgen2_A_I1068 (.Y(N2309), .A(N5636), .B(N5635), .S0(N5658));
MXI2XL addgen2_A_I1069 (.Y(N566), .A(N5660), .B(N5659), .S0(N2309));
MXI2XL addgen2_A_I1070 (.Y(N2318), .A(N5637), .B(N5636), .S0(N5658));
MXI2XL addgen2_A_I1071 (.Y(N567), .A(N5660), .B(N5659), .S0(N2318));
MXI2XL addgen2_A_I1072 (.Y(N2327), .A(N5638), .B(N5637), .S0(N5658));
MXI2XL addgen2_A_I1073 (.Y(N568), .A(N5660), .B(N5659), .S0(N2327));
MXI2XL addgen2_A_I1074 (.Y(N2336), .A(N5639), .B(N5638), .S0(N5658));
MXI2XL addgen2_A_I1075 (.Y(N569), .A(N5660), .B(N5659), .S0(N2336));
MXI2XL addgen2_A_I1076 (.Y(N2345), .A(N5640), .B(N5639), .S0(N5658));
MXI2XL addgen2_A_I1077 (.Y(N570), .A(N5660), .B(N5659), .S0(N2345));
MXI2XL addgen2_A_I1078 (.Y(N2354), .A(N5641), .B(N5640), .S0(N5658));
MXI2XL addgen2_A_I1079 (.Y(N571), .A(N5660), .B(N5659), .S0(N2354));
MXI2XL addgen2_A_I1080 (.Y(N2363), .A(N5642), .B(N5641), .S0(N5658));
MXI2XL addgen2_A_I1081 (.Y(N572), .A(N5660), .B(N5659), .S0(N2363));
MXI2XL addgen2_A_I1082 (.Y(N2372), .A(N5643), .B(N5642), .S0(N5658));
MXI2XL addgen2_A_I1083 (.Y(N573), .A(N5660), .B(N5659), .S0(N2372));
MXI2XL addgen2_A_I1084 (.Y(N2381), .A(N5644), .B(N5643), .S0(N5658));
MXI2XL addgen2_A_I1085 (.Y(N574), .A(N5660), .B(N5659), .S0(N2381));
MXI2XL addgen2_A_I1086 (.Y(N2390), .A(N5645), .B(N5644), .S0(N5658));
MXI2XL addgen2_A_I1087 (.Y(N575), .A(N5660), .B(N5659), .S0(N2390));
MXI2XL addgen2_A_I1088 (.Y(N2399), .A(N5646), .B(N5645), .S0(N5658));
MXI2XL addgen2_A_I1089 (.Y(N576), .A(N5660), .B(N5659), .S0(N2399));
MXI2XL addgen2_A_I1090 (.Y(N2408), .A(N5647), .B(N5646), .S0(N5658));
MXI2XL addgen2_A_I1091 (.Y(N577), .A(N5660), .B(N5659), .S0(N2408));
MXI2XL addgen2_A_I1092 (.Y(N2417), .A(N5648), .B(N5647), .S0(N5658));
MXI2XL addgen2_A_I1093 (.Y(N578), .A(N5660), .B(N5659), .S0(N2417));
MXI2XL addgen2_A_I1094 (.Y(N2426), .A(N5649), .B(N5648), .S0(N5658));
MXI2XL addgen2_A_I1095 (.Y(N579), .A(N5660), .B(N5659), .S0(N2426));
MXI2XL addgen2_A_I1096 (.Y(N2435), .A(N5650), .B(N5649), .S0(N5658));
MXI2XL addgen2_A_I1097 (.Y(N580), .A(N5660), .B(N5659), .S0(N2435));
MXI2XL addgen2_A_I1098 (.Y(N2444), .A(N5651), .B(N5650), .S0(N5658));
MXI2XL addgen2_A_I1099 (.Y(N581), .A(N5660), .B(N5659), .S0(N2444));
MXI2XL addgen2_A_I1100 (.Y(N2453), .A(N5652), .B(N5651), .S0(N5658));
MXI2XL addgen2_A_I1101 (.Y(N582), .A(N5660), .B(N5659), .S0(N2453));
MXI2XL addgen2_A_I1102 (.Y(N2462), .A(N5653), .B(N5652), .S0(N5658));
MXI2XL addgen2_A_I1103 (.Y(N583), .A(N5660), .B(N5659), .S0(N2462));
MXI2XL addgen2_A_I1104 (.Y(N2471), .A(N5654), .B(N5653), .S0(N5658));
MXI2XL addgen2_A_I1105 (.Y(N584), .A(N5660), .B(N5659), .S0(N2471));
NAND2XL addgen2_A_I1106 (.Y(N2480), .A(N5654), .B(N5658));
MXI2XL addgen2_A_I1107 (.Y(N585), .A(N5660), .B(N5659), .S0(N2480));
XNOR2X1 enc2_A_I1108 (.Y(N589), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
NOR2XL enc2_A_I1110 (.Y(N2491), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
OAI2BB1X1 enc2_A_I1825 (.Y(N588), .A0N(inst_cellmath__203_0_in1[20]), .A1N(inst_cellmath__203_0_in1[19]), .B0(inst_cellmath__203_0_in1[21]));
INVXL inst_cellmath__203_0_I1865 (.Y(N5661), .A(N588));
OR2XL inst_cellmath__203_0_I1969 (.Y(N5664), .A(N2491), .B(inst_cellmath__203_0_in1[21]));
INVXL inst_cellmath__203_0_I1869 (.Y(N5665), .A(N5661));
NOR2XL addgen2_A_I1113 (.Y(N2502), .A(N5635), .B(N589));
MXI2XL addgen2_A_I1114 (.Y(N595), .A(N5665), .B(N5664), .S0(N2502));
MXI2XL addgen2_A_I1115 (.Y(N2511), .A(N5636), .B(N5635), .S0(N589));
MXI2XL addgen2_A_I1116 (.Y(N596), .A(N5665), .B(N5664), .S0(N2511));
MXI2XL addgen2_A_I1117 (.Y(N2520), .A(N5637), .B(N5636), .S0(N589));
MXI2XL addgen2_A_I1118 (.Y(N597), .A(N5665), .B(N5664), .S0(N2520));
MXI2XL addgen2_A_I1119 (.Y(N2529), .A(N5638), .B(N5637), .S0(N589));
MXI2XL addgen2_A_I1120 (.Y(N598), .A(N5665), .B(N5664), .S0(N2529));
MXI2XL addgen2_A_I1121 (.Y(N2538), .A(N5639), .B(N5638), .S0(N589));
MXI2XL addgen2_A_I1122 (.Y(N599), .A(N5665), .B(N5664), .S0(N2538));
MXI2XL addgen2_A_I1123 (.Y(N2547), .A(N5640), .B(N5639), .S0(N589));
MXI2XL addgen2_A_I1124 (.Y(N600), .A(N5665), .B(N5664), .S0(N2547));
MXI2XL addgen2_A_I1125 (.Y(N2556), .A(N5641), .B(N5640), .S0(N589));
MXI2XL addgen2_A_I1126 (.Y(N601), .A(N5665), .B(N5664), .S0(N2556));
MXI2XL addgen2_A_I1127 (.Y(N2565), .A(N5642), .B(N5641), .S0(N589));
MXI2XL addgen2_A_I1128 (.Y(N602), .A(N5665), .B(N5664), .S0(N2565));
MXI2XL addgen2_A_I1129 (.Y(N2574), .A(N5643), .B(N5642), .S0(N589));
MXI2XL addgen2_A_I1130 (.Y(N603), .A(N5665), .B(N5664), .S0(N2574));
MXI2XL addgen2_A_I1131 (.Y(N2583), .A(N5644), .B(N5643), .S0(N589));
MXI2XL addgen2_A_I1132 (.Y(N604), .A(N5665), .B(N5664), .S0(N2583));
MXI2XL addgen2_A_I1133 (.Y(N2592), .A(N5645), .B(N5644), .S0(N589));
MXI2XL addgen2_A_I1134 (.Y(N605), .A(N5665), .B(N5664), .S0(N2592));
MXI2XL addgen2_A_I1135 (.Y(N2601), .A(N5646), .B(N5645), .S0(N589));
MXI2XL addgen2_A_I1136 (.Y(N606), .A(N5665), .B(N5664), .S0(N2601));
MXI2XL addgen2_A_I1137 (.Y(N2610), .A(N5647), .B(N5646), .S0(N589));
MXI2XL addgen2_A_I1138 (.Y(N607), .A(N5665), .B(N5664), .S0(N2610));
MXI2XL addgen2_A_I1139 (.Y(N2619), .A(N5648), .B(N5647), .S0(N589));
MXI2XL addgen2_A_I1140 (.Y(N608), .A(N5665), .B(N5664), .S0(N2619));
MXI2XL addgen2_A_I1141 (.Y(N2628), .A(N5649), .B(N5648), .S0(N589));
MXI2XL addgen2_A_I1142 (.Y(N609), .A(N5665), .B(N5664), .S0(N2628));
MXI2XL addgen2_A_I1143 (.Y(N2637), .A(N5650), .B(N5649), .S0(N589));
MXI2XL addgen2_A_I1144 (.Y(N610), .A(N5665), .B(N5664), .S0(N2637));
MXI2XL addgen2_A_I1145 (.Y(N2646), .A(N5651), .B(N5650), .S0(N589));
MXI2XL addgen2_A_I1146 (.Y(N611), .A(N5665), .B(N5664), .S0(N2646));
MXI2XL addgen2_A_I1147 (.Y(N2655), .A(N5652), .B(N5651), .S0(N589));
MXI2XL addgen2_A_I1148 (.Y(N612), .A(N5665), .B(N5664), .S0(N2655));
MXI2XL addgen2_A_I1149 (.Y(N2664), .A(N5653), .B(N5652), .S0(N589));
MXI2XL addgen2_A_I1150 (.Y(N613), .A(N5665), .B(N5664), .S0(N2664));
MXI2XL addgen2_A_I1151 (.Y(N2673), .A(N5654), .B(N5653), .S0(N589));
MXI2XL addgen2_A_I1152 (.Y(N614), .A(N5665), .B(N5664), .S0(N2673));
NAND2XL addgen2_A_I1153 (.Y(N2682), .A(N5654), .B(N589));
MXI2XL addgen2_A_I1154 (.Y(N615), .A(N5665), .B(N5664), .S0(N2682));
XNOR2X1 enc2_A_I1155 (.Y(N619), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
NOR2XL enc2_A_I1157 (.Y(N2693), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
OAI2BB1X1 enc2_A_I1826 (.Y(N618), .A0N(inst_cellmath__203_0_in1[22]), .A1N(inst_cellmath__203_0_in1[21]), .B0(inst_cellmath__203_0_in1[23]));
INVXL inst_cellmath__203_0_I1870 (.Y(N5666), .A(N618));
OR2XL inst_cellmath__203_0_I1970 (.Y(N5669), .A(N2693), .B(inst_cellmath__203_0_in1[23]));
INVXL inst_cellmath__203_0_I1874 (.Y(N5670), .A(N5666));
NOR2XL addgen2_A_I1160 (.Y(N2704), .A(N5635), .B(N619));
MXI2XL addgen2_A_I1161 (.Y(N625), .A(N5670), .B(N5669), .S0(N2704));
MXI2XL addgen2_A_I1162 (.Y(N2713), .A(N5636), .B(N5635), .S0(N619));
MXI2XL addgen2_A_I1163 (.Y(N626), .A(N5670), .B(N5669), .S0(N2713));
MXI2XL addgen2_A_I1164 (.Y(N2722), .A(N5637), .B(N5636), .S0(N619));
MXI2XL addgen2_A_I1165 (.Y(N627), .A(N5670), .B(N5669), .S0(N2722));
MXI2XL addgen2_A_I1166 (.Y(N2731), .A(N5638), .B(N5637), .S0(N619));
MXI2XL addgen2_A_I1167 (.Y(N628), .A(N5670), .B(N5669), .S0(N2731));
MXI2XL addgen2_A_I1168 (.Y(N2740), .A(N5639), .B(N5638), .S0(N619));
MXI2XL addgen2_A_I1169 (.Y(N629), .A(N5670), .B(N5669), .S0(N2740));
MXI2XL addgen2_A_I1170 (.Y(N2749), .A(N5640), .B(N5639), .S0(N619));
MXI2XL addgen2_A_I1171 (.Y(N630), .A(N5670), .B(N5669), .S0(N2749));
MXI2XL addgen2_A_I1172 (.Y(N2758), .A(N5641), .B(N5640), .S0(N619));
MXI2XL addgen2_A_I1173 (.Y(N631), .A(N5670), .B(N5669), .S0(N2758));
MXI2XL addgen2_A_I1174 (.Y(N2767), .A(N5642), .B(N5641), .S0(N619));
MXI2XL addgen2_A_I1175 (.Y(N632), .A(N5670), .B(N5669), .S0(N2767));
MXI2XL addgen2_A_I1176 (.Y(N2776), .A(N5643), .B(N5642), .S0(N619));
MXI2XL addgen2_A_I1177 (.Y(N633), .A(N5670), .B(N5669), .S0(N2776));
MXI2XL addgen2_A_I1178 (.Y(N2785), .A(N5644), .B(N5643), .S0(N619));
MXI2XL addgen2_A_I1179 (.Y(N634), .A(N5670), .B(N5669), .S0(N2785));
MXI2XL addgen2_A_I1180 (.Y(N2794), .A(N5645), .B(N5644), .S0(N619));
MXI2XL addgen2_A_I1181 (.Y(N635), .A(N5670), .B(N5669), .S0(N2794));
MXI2XL addgen2_A_I1182 (.Y(N2803), .A(N5646), .B(N5645), .S0(N619));
MXI2XL addgen2_A_I1183 (.Y(N636), .A(N5670), .B(N5669), .S0(N2803));
MXI2XL addgen2_A_I1184 (.Y(N2812), .A(N5647), .B(N5646), .S0(N619));
MXI2XL addgen2_A_I1185 (.Y(N637), .A(N5670), .B(N5669), .S0(N2812));
MXI2XL addgen2_A_I1186 (.Y(N2821), .A(N5648), .B(N5647), .S0(N619));
MXI2XL addgen2_A_I1187 (.Y(N638), .A(N5670), .B(N5669), .S0(N2821));
MXI2XL addgen2_A_I1188 (.Y(N2830), .A(N5649), .B(N5648), .S0(N619));
MXI2XL addgen2_A_I1189 (.Y(N639), .A(N5670), .B(N5669), .S0(N2830));
MXI2XL addgen2_A_I1190 (.Y(N2839), .A(N5650), .B(N5649), .S0(N619));
MXI2XL addgen2_A_I1191 (.Y(N640), .A(N5670), .B(N5669), .S0(N2839));
MXI2XL addgen2_A_I1192 (.Y(N2848), .A(N5651), .B(N5650), .S0(N619));
MXI2XL addgen2_A_I1193 (.Y(N641), .A(N5670), .B(N5669), .S0(N2848));
MXI2XL addgen2_A_I1194 (.Y(N2857), .A(N5652), .B(N5651), .S0(N619));
MXI2XL addgen2_A_I1195 (.Y(N642), .A(N5670), .B(N5669), .S0(N2857));
MXI2XL addgen2_A_I1196 (.Y(N2866), .A(N5653), .B(N5652), .S0(N619));
MXI2XL addgen2_A_I1197 (.Y(N643), .A(N5670), .B(N5669), .S0(N2866));
MXI2XL addgen2_A_I1198 (.Y(N2875), .A(N5654), .B(N5653), .S0(N619));
MXI2XL addgen2_A_I1199 (.Y(N644), .A(N5670), .B(N5669), .S0(N2875));
NAND2XL addgen2_A_I1200 (.Y(N2884), .A(N5654), .B(N619));
MXI2XL addgen2_A_I1201 (.Y(N645), .A(N5670), .B(N5669), .S0(N2884));
XNOR2X1 enc2_A_I1202 (.Y(N649), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
NOR2XL enc2_A_I1204 (.Y(N2895), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
OAI2BB1X1 enc2_A_I1827 (.Y(N648), .A0N(inst_cellmath__203_0_in1[24]), .A1N(inst_cellmath__203_0_in1[23]), .B0(inst_cellmath__203_0_in1[25]));
INVXL inst_cellmath__203_0_I1875 (.Y(N5671), .A(N648));
OR2XL inst_cellmath__203_0_I1971 (.Y(N5674), .A(N2895), .B(inst_cellmath__203_0_in1[25]));
INVXL inst_cellmath__203_0_I1879 (.Y(N5675), .A(N5671));
NOR2XL addgen2_A_I1207 (.Y(N2906), .A(N5635), .B(N649));
MXI2XL addgen2_A_I1208 (.Y(N655), .A(N5675), .B(N5674), .S0(N2906));
MXI2XL addgen2_A_I1209 (.Y(N2915), .A(N5636), .B(N5635), .S0(N649));
MXI2XL addgen2_A_I1210 (.Y(N656), .A(N5675), .B(N5674), .S0(N2915));
MXI2XL addgen2_A_I1211 (.Y(N2924), .A(N5637), .B(N5636), .S0(N649));
MXI2XL addgen2_A_I1212 (.Y(N657), .A(N5675), .B(N5674), .S0(N2924));
MXI2XL addgen2_A_I1213 (.Y(N2933), .A(N5638), .B(N5637), .S0(N649));
MXI2XL addgen2_A_I1214 (.Y(N658), .A(N5675), .B(N5674), .S0(N2933));
MXI2XL addgen2_A_I1215 (.Y(N2942), .A(N5639), .B(N5638), .S0(N649));
MXI2XL addgen2_A_I1216 (.Y(N659), .A(N5675), .B(N5674), .S0(N2942));
MXI2XL addgen2_A_I1217 (.Y(N2951), .A(N5640), .B(N5639), .S0(N649));
MXI2XL addgen2_A_I1218 (.Y(N660), .A(N5675), .B(N5674), .S0(N2951));
MXI2XL addgen2_A_I1219 (.Y(N2960), .A(N5641), .B(N5640), .S0(N649));
MXI2XL addgen2_A_I1220 (.Y(N661), .A(N5675), .B(N5674), .S0(N2960));
MXI2XL addgen2_A_I1221 (.Y(N2969), .A(N5642), .B(N5641), .S0(N649));
MXI2XL addgen2_A_I1222 (.Y(N662), .A(N5675), .B(N5674), .S0(N2969));
MXI2XL addgen2_A_I1223 (.Y(N2978), .A(N5643), .B(N5642), .S0(N649));
MXI2XL addgen2_A_I1224 (.Y(N663), .A(N5675), .B(N5674), .S0(N2978));
MXI2XL addgen2_A_I1225 (.Y(N2987), .A(N5644), .B(N5643), .S0(N649));
MXI2XL addgen2_A_I1226 (.Y(N664), .A(N5675), .B(N5674), .S0(N2987));
MXI2XL addgen2_A_I1227 (.Y(N2996), .A(N5645), .B(N5644), .S0(N649));
MXI2XL addgen2_A_I1228 (.Y(N665), .A(N5675), .B(N5674), .S0(N2996));
MXI2XL addgen2_A_I1229 (.Y(N3005), .A(N5646), .B(N5645), .S0(N649));
MXI2XL addgen2_A_I1230 (.Y(N666), .A(N5675), .B(N5674), .S0(N3005));
MXI2XL addgen2_A_I1231 (.Y(N3014), .A(N5647), .B(N5646), .S0(N649));
MXI2XL addgen2_A_I1232 (.Y(N667), .A(N5675), .B(N5674), .S0(N3014));
MXI2XL addgen2_A_I1233 (.Y(N3023), .A(N5648), .B(N5647), .S0(N649));
MXI2XL addgen2_A_I1234 (.Y(N668), .A(N5675), .B(N5674), .S0(N3023));
MXI2XL addgen2_A_I1235 (.Y(N3032), .A(N5649), .B(N5648), .S0(N649));
MXI2XL addgen2_A_I1236 (.Y(N669), .A(N5675), .B(N5674), .S0(N3032));
MXI2XL addgen2_A_I1237 (.Y(N3041), .A(N5650), .B(N5649), .S0(N649));
MXI2XL addgen2_A_I1238 (.Y(N670), .A(N5675), .B(N5674), .S0(N3041));
MXI2XL addgen2_A_I1239 (.Y(N3050), .A(N5651), .B(N5650), .S0(N649));
MXI2XL addgen2_A_I1240 (.Y(N671), .A(N5675), .B(N5674), .S0(N3050));
MXI2XL addgen2_A_I1241 (.Y(N3059), .A(N5652), .B(N5651), .S0(N649));
MXI2XL addgen2_A_I1242 (.Y(N672), .A(N5675), .B(N5674), .S0(N3059));
MXI2XL addgen2_A_I1243 (.Y(N3068), .A(N5653), .B(N5652), .S0(N649));
MXI2XL addgen2_A_I1244 (.Y(N673), .A(N5675), .B(N5674), .S0(N3068));
MXI2XL addgen2_A_I1245 (.Y(N3077), .A(N5654), .B(N5653), .S0(N649));
MXI2XL addgen2_A_I1246 (.Y(N674), .A(N5675), .B(N5674), .S0(N3077));
NAND2XL addgen2_A_I1247 (.Y(N3086), .A(N5654), .B(N649));
MXI2XL addgen2_A_I1248 (.Y(N675), .A(N5675), .B(N5674), .S0(N3086));
XNOR2X1 enc2_A_I1249 (.Y(N679), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
NOR2XL enc2_A_I1251 (.Y(N3097), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
OAI2BB1X1 enc2_A_I1828 (.Y(N678), .A0N(inst_cellmath__203_0_in1[26]), .A1N(inst_cellmath__203_0_in1[25]), .B0(inst_cellmath__203_0_in1[27]));
INVXL inst_cellmath__203_0_I1880 (.Y(N5676), .A(N678));
OR2XL inst_cellmath__203_0_I1972 (.Y(N5679), .A(N3097), .B(inst_cellmath__203_0_in1[27]));
INVXL inst_cellmath__203_0_I1884 (.Y(N5680), .A(N5676));
NOR2XL addgen2_A_I1254 (.Y(N3108), .A(N5635), .B(N679));
MXI2XL addgen2_A_I1255 (.Y(N685), .A(N5680), .B(N5679), .S0(N3108));
MXI2XL addgen2_A_I1256 (.Y(N3117), .A(N5636), .B(N5635), .S0(N679));
MXI2XL addgen2_A_I1257 (.Y(N686), .A(N5680), .B(N5679), .S0(N3117));
MXI2XL addgen2_A_I1258 (.Y(N3126), .A(N5637), .B(N5636), .S0(N679));
MXI2XL addgen2_A_I1259 (.Y(N687), .A(N5680), .B(N5679), .S0(N3126));
MXI2XL addgen2_A_I1260 (.Y(N3135), .A(N5638), .B(N5637), .S0(N679));
MXI2XL addgen2_A_I1261 (.Y(N688), .A(N5680), .B(N5679), .S0(N3135));
MXI2XL addgen2_A_I1262 (.Y(N3144), .A(N5639), .B(N5638), .S0(N679));
MXI2XL addgen2_A_I1263 (.Y(N689), .A(N5680), .B(N5679), .S0(N3144));
MXI2XL addgen2_A_I1264 (.Y(N3153), .A(N5640), .B(N5639), .S0(N679));
MXI2XL addgen2_A_I1265 (.Y(N690), .A(N5680), .B(N5679), .S0(N3153));
MXI2XL addgen2_A_I1266 (.Y(N3162), .A(N5641), .B(N5640), .S0(N679));
MXI2XL addgen2_A_I1267 (.Y(N691), .A(N5680), .B(N5679), .S0(N3162));
MXI2XL addgen2_A_I1268 (.Y(N3171), .A(N5642), .B(N5641), .S0(N679));
MXI2XL addgen2_A_I1269 (.Y(N692), .A(N5680), .B(N5679), .S0(N3171));
MXI2XL addgen2_A_I1270 (.Y(N3180), .A(N5643), .B(N5642), .S0(N679));
MXI2XL addgen2_A_I1271 (.Y(N693), .A(N5680), .B(N5679), .S0(N3180));
MXI2XL addgen2_A_I1272 (.Y(N3189), .A(N5644), .B(N5643), .S0(N679));
MXI2XL addgen2_A_I1273 (.Y(N694), .A(N5680), .B(N5679), .S0(N3189));
MXI2XL addgen2_A_I1274 (.Y(N3198), .A(N5645), .B(N5644), .S0(N679));
MXI2XL addgen2_A_I1275 (.Y(N695), .A(N5680), .B(N5679), .S0(N3198));
MXI2XL addgen2_A_I1276 (.Y(N3207), .A(N5646), .B(N5645), .S0(N679));
MXI2XL addgen2_A_I1277 (.Y(N696), .A(N5680), .B(N5679), .S0(N3207));
MXI2XL addgen2_A_I1278 (.Y(N3216), .A(N5647), .B(N5646), .S0(N679));
MXI2XL addgen2_A_I1279 (.Y(N697), .A(N5680), .B(N5679), .S0(N3216));
MXI2XL addgen2_A_I1280 (.Y(N3225), .A(N5648), .B(N5647), .S0(N679));
MXI2XL addgen2_A_I1281 (.Y(N698), .A(N5680), .B(N5679), .S0(N3225));
MXI2XL addgen2_A_I1282 (.Y(N3234), .A(N5649), .B(N5648), .S0(N679));
MXI2XL addgen2_A_I1283 (.Y(N699), .A(N5680), .B(N5679), .S0(N3234));
MXI2XL addgen2_A_I1284 (.Y(N3243), .A(N5650), .B(N5649), .S0(N679));
MXI2XL addgen2_A_I1285 (.Y(N700), .A(N5680), .B(N5679), .S0(N3243));
MXI2XL addgen2_A_I1286 (.Y(N3252), .A(N5651), .B(N5650), .S0(N679));
MXI2XL addgen2_A_I1287 (.Y(N701), .A(N5680), .B(N5679), .S0(N3252));
MXI2XL addgen2_A_I1288 (.Y(N3261), .A(N5652), .B(N5651), .S0(N679));
MXI2XL addgen2_A_I1289 (.Y(N702), .A(N5680), .B(N5679), .S0(N3261));
MXI2XL addgen2_A_I1290 (.Y(N3270), .A(N5653), .B(N5652), .S0(N679));
MXI2XL addgen2_A_I1291 (.Y(N703), .A(N5680), .B(N5679), .S0(N3270));
MXI2XL addgen2_A_I1292 (.Y(N3279), .A(N5654), .B(N5653), .S0(N679));
MXI2XL addgen2_A_I1293 (.Y(N704), .A(N5680), .B(N5679), .S0(N3279));
NAND2XL addgen2_A_I1294 (.Y(N3288), .A(N5654), .B(N679));
MXI2XL addgen2_A_I1295 (.Y(N705), .A(N5680), .B(N5679), .S0(N3288));
XNOR2X1 enc2_A_I1296 (.Y(N709), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
NOR2XL enc2_A_I1298 (.Y(N3299), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
OAI2BB1X1 enc2_A_I1829 (.Y(N708), .A0N(inst_cellmath__203_0_in1[28]), .A1N(inst_cellmath__203_0_in1[27]), .B0(inst_cellmath__203_0_in1[29]));
INVXL inst_cellmath__203_0_I1885 (.Y(N5681), .A(N708));
OR2XL inst_cellmath__203_0_I1973 (.Y(N5684), .A(N3299), .B(inst_cellmath__203_0_in1[29]));
INVXL inst_cellmath__203_0_I1889 (.Y(N5685), .A(N5681));
NOR2XL addgen2_A_I1301 (.Y(N3310), .A(N5635), .B(N709));
MXI2XL addgen2_A_I1302 (.Y(N715), .A(N5685), .B(N5684), .S0(N3310));
MXI2XL addgen2_A_I1303 (.Y(N3319), .A(N5636), .B(N5635), .S0(N709));
MXI2XL addgen2_A_I1304 (.Y(N716), .A(N5685), .B(N5684), .S0(N3319));
MXI2XL addgen2_A_I1305 (.Y(N3328), .A(N5637), .B(N5636), .S0(N709));
MXI2XL addgen2_A_I1306 (.Y(N717), .A(N5685), .B(N5684), .S0(N3328));
MXI2XL addgen2_A_I1307 (.Y(N3337), .A(N5638), .B(N5637), .S0(N709));
MXI2XL addgen2_A_I1308 (.Y(N718), .A(N5685), .B(N5684), .S0(N3337));
MXI2XL addgen2_A_I1309 (.Y(N3346), .A(N5639), .B(N5638), .S0(N709));
MXI2XL addgen2_A_I1310 (.Y(N719), .A(N5685), .B(N5684), .S0(N3346));
MXI2XL addgen2_A_I1311 (.Y(N3355), .A(N5640), .B(N5639), .S0(N709));
MXI2XL addgen2_A_I1312 (.Y(N720), .A(N5685), .B(N5684), .S0(N3355));
MXI2XL addgen2_A_I1313 (.Y(N3364), .A(N5641), .B(N5640), .S0(N709));
MXI2XL addgen2_A_I1314 (.Y(N721), .A(N5685), .B(N5684), .S0(N3364));
MXI2XL addgen2_A_I1315 (.Y(N3373), .A(N5642), .B(N5641), .S0(N709));
MXI2XL addgen2_A_I1316 (.Y(N722), .A(N5685), .B(N5684), .S0(N3373));
MXI2XL addgen2_A_I1317 (.Y(N3382), .A(N5643), .B(N5642), .S0(N709));
MXI2XL addgen2_A_I1318 (.Y(N723), .A(N5685), .B(N5684), .S0(N3382));
MXI2XL addgen2_A_I1319 (.Y(N3391), .A(N5644), .B(N5643), .S0(N709));
MXI2XL addgen2_A_I1320 (.Y(N724), .A(N5685), .B(N5684), .S0(N3391));
MXI2XL addgen2_A_I1321 (.Y(N3400), .A(N5645), .B(N5644), .S0(N709));
MXI2XL addgen2_A_I1322 (.Y(N725), .A(N5685), .B(N5684), .S0(N3400));
MXI2XL addgen2_A_I1323 (.Y(N3409), .A(N5646), .B(N5645), .S0(N709));
MXI2XL addgen2_A_I1324 (.Y(N726), .A(N5685), .B(N5684), .S0(N3409));
MXI2XL addgen2_A_I1325 (.Y(N3418), .A(N5647), .B(N5646), .S0(N709));
MXI2XL addgen2_A_I1326 (.Y(N727), .A(N5685), .B(N5684), .S0(N3418));
MXI2XL addgen2_A_I1327 (.Y(N3427), .A(N5648), .B(N5647), .S0(N709));
MXI2XL addgen2_A_I1328 (.Y(N728), .A(N5685), .B(N5684), .S0(N3427));
MXI2XL addgen2_A_I1329 (.Y(N3436), .A(N5649), .B(N5648), .S0(N709));
MXI2XL addgen2_A_I1330 (.Y(N729), .A(N5685), .B(N5684), .S0(N3436));
MXI2XL addgen2_A_I1331 (.Y(N3445), .A(N5650), .B(N5649), .S0(N709));
MXI2XL addgen2_A_I1332 (.Y(N730), .A(N5685), .B(N5684), .S0(N3445));
MXI2XL addgen2_A_I1333 (.Y(N3454), .A(N5651), .B(N5650), .S0(N709));
MXI2XL addgen2_A_I1334 (.Y(N731), .A(N5685), .B(N5684), .S0(N3454));
MXI2XL addgen2_A_I1335 (.Y(N3463), .A(N5652), .B(N5651), .S0(N709));
MXI2XL addgen2_A_I1336 (.Y(N732), .A(N5685), .B(N5684), .S0(N3463));
MXI2XL addgen2_A_I1337 (.Y(N3472), .A(N5653), .B(N5652), .S0(N709));
MXI2XL addgen2_A_I1338 (.Y(N733), .A(N5685), .B(N5684), .S0(N3472));
MXI2XL addgen2_A_I1339 (.Y(N3481), .A(N5654), .B(N5653), .S0(N709));
MXI2XL addgen2_A_I1340 (.Y(N734), .A(N5685), .B(N5684), .S0(N3481));
NAND2XL addgen2_A_I1341 (.Y(N3490), .A(N5654), .B(N709));
MXI2XL addgen2_A_I1342 (.Y(N735), .A(N5685), .B(N5684), .S0(N3490));
XNOR2X1 enc2_A_I1343 (.Y(N739), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
NOR2XL enc2_A_I1345 (.Y(N3501), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
OAI2BB1X1 enc2_A_I1830 (.Y(N738), .A0N(inst_cellmath__203_0_in1[30]), .A1N(inst_cellmath__203_0_in1[29]), .B0(inst_cellmath__203_0_in1[31]));
INVXL inst_cellmath__203_0_I1890 (.Y(N5686), .A(N738));
OR2XL inst_cellmath__203_0_I1974 (.Y(N5689), .A(N3501), .B(inst_cellmath__203_0_in1[31]));
INVXL inst_cellmath__203_0_I1894 (.Y(N5690), .A(N5686));
NOR2XL addgen2_A_I1348 (.Y(N3512), .A(N5635), .B(N739));
MXI2XL addgen2_A_I1349 (.Y(N745), .A(N5690), .B(N5689), .S0(N3512));
MXI2XL addgen2_A_I1350 (.Y(N3521), .A(N5636), .B(N5635), .S0(N739));
MXI2XL addgen2_A_I1351 (.Y(N746), .A(N5690), .B(N5689), .S0(N3521));
MXI2XL addgen2_A_I1352 (.Y(N3530), .A(N5637), .B(N5636), .S0(N739));
MXI2XL addgen2_A_I1353 (.Y(N747), .A(N5690), .B(N5689), .S0(N3530));
MXI2XL addgen2_A_I1354 (.Y(N3539), .A(N5638), .B(N5637), .S0(N739));
MXI2XL addgen2_A_I1355 (.Y(N748), .A(N5690), .B(N5689), .S0(N3539));
MXI2XL addgen2_A_I1356 (.Y(N3548), .A(N5639), .B(N5638), .S0(N739));
MXI2XL addgen2_A_I1357 (.Y(N749), .A(N5690), .B(N5689), .S0(N3548));
MXI2XL addgen2_A_I1358 (.Y(N3557), .A(N5640), .B(N5639), .S0(N739));
MXI2XL addgen2_A_I1359 (.Y(N750), .A(N5690), .B(N5689), .S0(N3557));
MXI2XL addgen2_A_I1360 (.Y(N3566), .A(N5641), .B(N5640), .S0(N739));
MXI2XL addgen2_A_I1361 (.Y(N751), .A(N5690), .B(N5689), .S0(N3566));
MXI2XL addgen2_A_I1362 (.Y(N3575), .A(N5642), .B(N5641), .S0(N739));
MXI2XL addgen2_A_I1363 (.Y(N752), .A(N5690), .B(N5689), .S0(N3575));
MXI2XL addgen2_A_I1364 (.Y(N3584), .A(N5643), .B(N5642), .S0(N739));
MXI2XL addgen2_A_I1365 (.Y(N753), .A(N5690), .B(N5689), .S0(N3584));
MXI2XL addgen2_A_I1366 (.Y(N3593), .A(N5644), .B(N5643), .S0(N739));
MXI2XL addgen2_A_I1367 (.Y(N754), .A(N5690), .B(N5689), .S0(N3593));
MXI2XL addgen2_A_I1368 (.Y(N3602), .A(N5645), .B(N5644), .S0(N739));
MXI2XL addgen2_A_I1369 (.Y(N755), .A(N5690), .B(N5689), .S0(N3602));
MXI2XL addgen2_A_I1370 (.Y(N3611), .A(N5646), .B(N5645), .S0(N739));
MXI2XL addgen2_A_I1371 (.Y(N756), .A(N5690), .B(N5689), .S0(N3611));
MXI2XL addgen2_A_I1372 (.Y(N3620), .A(N5647), .B(N5646), .S0(N739));
MXI2XL addgen2_A_I1373 (.Y(N757), .A(N5690), .B(N5689), .S0(N3620));
MXI2XL addgen2_A_I1374 (.Y(N3629), .A(N5648), .B(N5647), .S0(N739));
MXI2XL addgen2_A_I1375 (.Y(N758), .A(N5690), .B(N5689), .S0(N3629));
MXI2XL addgen2_A_I1376 (.Y(N3638), .A(N5649), .B(N5648), .S0(N739));
MXI2XL addgen2_A_I1377 (.Y(N759), .A(N5690), .B(N5689), .S0(N3638));
MXI2XL addgen2_A_I1378 (.Y(N3647), .A(N5650), .B(N5649), .S0(N739));
MXI2XL addgen2_A_I1379 (.Y(N760), .A(N5690), .B(N5689), .S0(N3647));
MXI2XL addgen2_A_I1380 (.Y(N3656), .A(N5651), .B(N5650), .S0(N739));
MXI2XL addgen2_A_I1381 (.Y(N761), .A(N5690), .B(N5689), .S0(N3656));
MXI2XL addgen2_A_I1382 (.Y(N3665), .A(N5652), .B(N5651), .S0(N739));
MXI2XL addgen2_A_I1383 (.Y(N762), .A(N5690), .B(N5689), .S0(N3665));
MXI2XL addgen2_A_I1384 (.Y(N3674), .A(N5653), .B(N5652), .S0(N739));
MXI2XL addgen2_A_I1385 (.Y(N763), .A(N5690), .B(N5689), .S0(N3674));
MXI2XL addgen2_A_I1386 (.Y(N3683), .A(N5654), .B(N5653), .S0(N739));
MXI2XL addgen2_A_I1387 (.Y(N764), .A(N5690), .B(N5689), .S0(N3683));
NAND2XL addgen2_A_I1388 (.Y(N3692), .A(N5654), .B(N739));
MXI2XL addgen2_A_I1389 (.Y(N765), .A(N5690), .B(N5689), .S0(N3692));
ADDHX1 inst_cellmath__203_0_I281 (.CO(N770), .S(N768), .A(inst_cellmath__203_0_in1[32]), .B(inst_cellmath__203_0_in1[31]));
INVXL inst_cellmath__203_0_I1895 (.Y(N5691), .A(N768));
INVXL inst_cellmath__203_0_I1896 (.Y(N5692), .A(N770));
NOR2XL inst_cellmath__203_0_I285 (.Y(N779), .A(N5691), .B(N5635));
OAI22XL inst_cellmath__203_0_I286 (.Y(N781), .A0(N5635), .A1(N5692), .B0(N5691), .B1(N5636));
OAI22XL inst_cellmath__203_0_I287 (.Y(N783), .A0(N5636), .A1(N5692), .B0(N5691), .B1(N5637));
OAI22XL inst_cellmath__203_0_I288 (.Y(N785), .A0(N5637), .A1(N5692), .B0(N5691), .B1(N5638));
OAI22XL inst_cellmath__203_0_I289 (.Y(N787), .A0(N5638), .A1(N5692), .B0(N5691), .B1(N5639));
OAI22XL inst_cellmath__203_0_I290 (.Y(N789), .A0(N5639), .A1(N5692), .B0(N5691), .B1(N5640));
OAI22XL inst_cellmath__203_0_I291 (.Y(N791), .A0(N5640), .A1(N5692), .B0(N5691), .B1(N5641));
OAI22XL inst_cellmath__203_0_I292 (.Y(N793), .A0(N5641), .A1(N5692), .B0(N5691), .B1(N5642));
OAI22XL inst_cellmath__203_0_I293 (.Y(N795), .A0(N5642), .A1(N5692), .B0(N5691), .B1(N5643));
OAI22XL inst_cellmath__203_0_I294 (.Y(N797), .A0(N5643), .A1(N5692), .B0(N5691), .B1(N5644));
OAI22XL inst_cellmath__203_0_I295 (.Y(N799), .A0(N5644), .A1(N5692), .B0(N5691), .B1(N5645));
OAI22XL inst_cellmath__203_0_I296 (.Y(N801), .A0(N5645), .A1(N5692), .B0(N5691), .B1(N5646));
OAI22XL inst_cellmath__203_0_I297 (.Y(N803), .A0(N5646), .A1(N5692), .B0(N5691), .B1(N5647));
OAI22XL inst_cellmath__203_0_I298 (.Y(N805), .A0(N5647), .A1(N5692), .B0(N5691), .B1(N5648));
OAI22XL inst_cellmath__203_0_I299 (.Y(N807), .A0(N5648), .A1(N5692), .B0(N5691), .B1(N5649));
OAI22XL inst_cellmath__203_0_I300 (.Y(N809), .A0(N5649), .A1(N5692), .B0(N5691), .B1(N5650));
OAI22XL inst_cellmath__203_0_I301 (.Y(N811), .A0(N5650), .A1(N5692), .B0(N5691), .B1(N5651));
OAI22XL inst_cellmath__203_0_I302 (.Y(N813), .A0(N5651), .A1(N5692), .B0(N5691), .B1(N5652));
OAI22XL inst_cellmath__203_0_I303 (.Y(N815), .A0(N5652), .A1(N5692), .B0(N5691), .B1(N5653));
OAI22XL inst_cellmath__203_0_I304 (.Y(N817), .A0(N5653), .A1(N5692), .B0(N5691), .B1(N5654));
OAI21XL inst_cellmath__203_0_I305 (.Y(N819), .A0(N5692), .A1(N5654), .B0(N5691));
AND2XL inst_cellmath__203_0_I306 (.Y(N1366), .A(N5692), .B(N5691));
INVXL inst_cellmath__203_0_I1897 (.Y(N5693), .A(inst_cellmath__203_0_in3[0]));
INVXL inst_cellmath__203_0_I1898 (.Y(N5694), .A(inst_cellmath__203_0_in3[1]));
INVXL inst_cellmath__203_0_I1899 (.Y(N5695), .A(inst_cellmath__203_0_in3[2]));
INVXL inst_cellmath__203_0_I1900 (.Y(N5696), .A(inst_cellmath__203_0_in3[3]));
INVXL inst_cellmath__203_0_I1901 (.Y(N5697), .A(inst_cellmath__203_0_in3[4]));
INVXL inst_cellmath__203_0_I1902 (.Y(N5698), .A(inst_cellmath__203_0_in3[5]));
INVXL inst_cellmath__203_0_I1903 (.Y(N5699), .A(inst_cellmath__203_0_in3[6]));
INVXL inst_cellmath__203_0_I1904 (.Y(N5700), .A(inst_cellmath__203_0_in3[7]));
INVXL inst_cellmath__203_0_I1905 (.Y(N5701), .A(inst_cellmath__203_0_in3[8]));
INVXL inst_cellmath__203_0_I1906 (.Y(N5702), .A(inst_cellmath__203_0_in3[9]));
INVXL inst_cellmath__203_0_I1907 (.Y(N5703), .A(inst_cellmath__203_0_in3[10]));
INVXL inst_cellmath__203_0_I1908 (.Y(N5704), .A(inst_cellmath__203_0_in3[11]));
INVXL inst_cellmath__203_0_I1909 (.Y(N5705), .A(inst_cellmath__203_0_in3[12]));
INVXL inst_cellmath__203_0_I1910 (.Y(N5706), .A(inst_cellmath__203_0_in3[13]));
INVXL inst_cellmath__203_0_I1911 (.Y(N5707), .A(inst_cellmath__203_0_in3[14]));
INVXL inst_cellmath__203_0_I1912 (.Y(N5708), .A(inst_cellmath__203_0_in3[15]));
INVXL inst_cellmath__203_0_I1913 (.Y(N5709), .A(inst_cellmath__203_0_in3[16]));
INVXL inst_cellmath__203_0_I1914 (.Y(N5710), .A(inst_cellmath__203_0_in3[17]));
INVXL inst_cellmath__203_0_I1915 (.Y(N5711), .A(inst_cellmath__203_0_in3[18]));
INVXL inst_cellmath__203_0_I1916 (.Y(N5712), .A(inst_cellmath__203_0_in3[19]));
INVXL inst_cellmath__203_0_I1917 (.Y(N5713), .A(inst_cellmath__203_0_in3[20]));
INVXL inst_cellmath__203_0_I1918 (.Y(N5714), .A(inst_cellmath__203_0_in3[21]));
INVXL inst_cellmath__203_0_I1919 (.Y(N5715), .A(inst_cellmath__203_0_in0[0]));
NOR2XL inst_cellmath__203_0_I382 (.Y(N1025), .A(N5715), .B(N5693));
NOR2XL inst_cellmath__203_0_I383 (.Y(N1027), .A(N5715), .B(N5694));
NOR2XL inst_cellmath__203_0_I384 (.Y(N1029), .A(N5715), .B(N5695));
NOR2XL inst_cellmath__203_0_I385 (.Y(N1031), .A(N5715), .B(N5696));
NOR2XL inst_cellmath__203_0_I386 (.Y(N1033), .A(N5715), .B(N5697));
NOR2XL inst_cellmath__203_0_I387 (.Y(N1035), .A(N5715), .B(N5698));
NOR2XL inst_cellmath__203_0_I388 (.Y(N1037), .A(N5715), .B(N5699));
NOR2XL inst_cellmath__203_0_I389 (.Y(N1039), .A(N5715), .B(N5700));
NOR2XL inst_cellmath__203_0_I390 (.Y(N1041), .A(N5715), .B(N5701));
NOR2XL inst_cellmath__203_0_I391 (.Y(N1043), .A(N5715), .B(N5702));
NOR2XL inst_cellmath__203_0_I392 (.Y(N1045), .A(N5715), .B(N5703));
NOR2XL inst_cellmath__203_0_I393 (.Y(N1047), .A(N5715), .B(N5704));
NOR2XL inst_cellmath__203_0_I394 (.Y(N1049), .A(N5715), .B(N5705));
NOR2XL inst_cellmath__203_0_I395 (.Y(N1051), .A(N5715), .B(N5706));
NOR2XL inst_cellmath__203_0_I396 (.Y(N1053), .A(N5715), .B(N5707));
NOR2XL inst_cellmath__203_0_I397 (.Y(N1055), .A(N5715), .B(N5708));
NOR2XL inst_cellmath__203_0_I398 (.Y(N1732), .A(N5715), .B(N5709));
NOR2XL inst_cellmath__203_0_I399 (.Y(N1059), .A(N5715), .B(N5710));
NOR2XL inst_cellmath__203_0_I400 (.Y(N1061), .A(N5715), .B(N5711));
NOR2XL inst_cellmath__203_0_I401 (.Y(N1798), .A(N5715), .B(N5712));
NOR2XL inst_cellmath__203_0_I402 (.Y(N1830), .A(N5715), .B(N5713));
NOR2XL inst_cellmath__203_0_I403 (.Y(N1067), .A(N5715), .B(N5714));
INVXL inst_cellmath__203_0_I1922 (.Y(N5718), .A(inst_cellmath__203_0_in0[1]));
NAND2BX1 inst_cellmath__203_0_I1975 (.Y(N5719), .AN(inst_cellmath__203_0_in0[2]), .B(inst_cellmath__203_0_in0[1]));
INVXL inst_cellmath__203_0_I1924 (.Y(N5720), .A(inst_cellmath__203_0_in0[2]));
NOR2XL addgen2_A_I1395 (.Y(N3714), .A(N5693), .B(N5718));
MXI2XL addgen2_A_I1396 (.Y(N1077), .A(N5720), .B(N5719), .S0(N3714));
MXI2XL addgen2_A_I1397 (.Y(N3723), .A(N5694), .B(N5693), .S0(N5718));
MXI2XL addgen2_A_I1398 (.Y(N1078), .A(N5720), .B(N5719), .S0(N3723));
MXI2XL addgen2_A_I1399 (.Y(N3732), .A(N5695), .B(N5694), .S0(N5718));
MXI2XL addgen2_A_I1400 (.Y(N1079), .A(N5720), .B(N5719), .S0(N3732));
MXI2XL addgen2_A_I1401 (.Y(N3741), .A(N5696), .B(N5695), .S0(N5718));
MXI2XL addgen2_A_I1402 (.Y(N1080), .A(N5720), .B(N5719), .S0(N3741));
MXI2XL addgen2_A_I1403 (.Y(N3750), .A(N5697), .B(N5696), .S0(N5718));
MXI2XL addgen2_A_I1404 (.Y(N1081), .A(N5720), .B(N5719), .S0(N3750));
MXI2XL addgen2_A_I1405 (.Y(N3759), .A(N5698), .B(N5697), .S0(N5718));
MXI2XL addgen2_A_I1406 (.Y(N1082), .A(N5720), .B(N5719), .S0(N3759));
MXI2XL addgen2_A_I1407 (.Y(N3768), .A(N5699), .B(N5698), .S0(N5718));
MXI2XL addgen2_A_I1408 (.Y(N1083), .A(N5720), .B(N5719), .S0(N3768));
MXI2XL addgen2_A_I1409 (.Y(N3777), .A(N5700), .B(N5699), .S0(N5718));
MXI2XL addgen2_A_I1410 (.Y(N1084), .A(N5720), .B(N5719), .S0(N3777));
MXI2XL addgen2_A_I1411 (.Y(N3786), .A(N5701), .B(N5700), .S0(N5718));
MXI2XL addgen2_A_I1412 (.Y(N1085), .A(N5720), .B(N5719), .S0(N3786));
MXI2XL addgen2_A_I1413 (.Y(N3795), .A(N5702), .B(N5701), .S0(N5718));
MXI2XL addgen2_A_I1414 (.Y(N1086), .A(N5720), .B(N5719), .S0(N3795));
MXI2XL addgen2_A_I1415 (.Y(N3804), .A(N5703), .B(N5702), .S0(N5718));
MXI2XL addgen2_A_I1416 (.Y(N1087), .A(N5720), .B(N5719), .S0(N3804));
MXI2XL addgen2_A_I1417 (.Y(N3813), .A(N5704), .B(N5703), .S0(N5718));
MXI2XL addgen2_A_I1418 (.Y(N1088), .A(N5720), .B(N5719), .S0(N3813));
MXI2XL addgen2_A_I1419 (.Y(N3822), .A(N5705), .B(N5704), .S0(N5718));
MXI2XL addgen2_A_I1420 (.Y(N1089), .A(N5720), .B(N5719), .S0(N3822));
MXI2XL addgen2_A_I1421 (.Y(N3831), .A(N5706), .B(N5705), .S0(N5718));
MXI2XL addgen2_A_I1422 (.Y(N1090), .A(N5720), .B(N5719), .S0(N3831));
MXI2XL addgen2_A_I1423 (.Y(N3840), .A(N5707), .B(N5706), .S0(N5718));
MXI2XL addgen2_A_I1424 (.Y(N1091), .A(N5720), .B(N5719), .S0(N3840));
MXI2XL addgen2_A_I1425 (.Y(N3849), .A(N5708), .B(N5707), .S0(N5718));
MXI2XL addgen2_A_I1426 (.Y(N1092), .A(N5720), .B(N5719), .S0(N3849));
MXI2XL addgen2_A_I1427 (.Y(N3858), .A(N5709), .B(N5708), .S0(N5718));
MXI2XL addgen2_A_I1428 (.Y(N1093), .A(N5720), .B(N5719), .S0(N3858));
MXI2XL addgen2_A_I1429 (.Y(N3867), .A(N5710), .B(N5709), .S0(N5718));
MXI2XL addgen2_A_I1430 (.Y(N1094), .A(N5720), .B(N5719), .S0(N3867));
MXI2XL addgen2_A_I1431 (.Y(N3876), .A(N5711), .B(N5710), .S0(N5718));
MXI2XL addgen2_A_I1432 (.Y(N1095), .A(N5720), .B(N5719), .S0(N3876));
MXI2XL addgen2_A_I1433 (.Y(N3885), .A(N5712), .B(N5711), .S0(N5718));
MXI2XL addgen2_A_I1434 (.Y(N1096), .A(N5720), .B(N5719), .S0(N3885));
MXI2XL addgen2_A_I1435 (.Y(N3894), .A(N5713), .B(N5712), .S0(N5718));
MXI2XL addgen2_A_I1436 (.Y(N1097), .A(N5720), .B(N5719), .S0(N3894));
MXI2XL addgen2_A_I1437 (.Y(N3903), .A(N5714), .B(N5713), .S0(N5718));
MXI2XL addgen2_A_I1438 (.Y(N1098), .A(N5720), .B(N5719), .S0(N3903));
NOR2BX1 addgen2_A_I1439 (.Y(N3912), .AN(N5718), .B(N5714));
MXI2XL addgen2_A_I1440 (.Y(N1099), .A(N5720), .B(N5719), .S0(N3912));
XNOR2X1 enc2_A_I1441 (.Y(N1103), .A(inst_cellmath__203_0_in0[3]), .B(inst_cellmath__203_0_in0[2]));
NOR2XL enc2_A_I1443 (.Y(N3923), .A(inst_cellmath__203_0_in0[3]), .B(inst_cellmath__203_0_in0[2]));
OAI2BB1X1 enc2_A_I1832 (.Y(N1102), .A0N(inst_cellmath__203_0_in0[3]), .A1N(inst_cellmath__203_0_in0[2]), .B0(inst_cellmath__203_0_in0[4]));
INVXL inst_cellmath__203_0_I1925 (.Y(N5721), .A(N1102));
OR2XL inst_cellmath__203_0_I1976 (.Y(N5724), .A(N3923), .B(inst_cellmath__203_0_in0[4]));
INVXL inst_cellmath__203_0_I1929 (.Y(N5725), .A(N5721));
NOR2XL addgen2_A_I1446 (.Y(N3934), .A(N5693), .B(N1103));
MXI2XL addgen2_A_I1447 (.Y(N1109), .A(N5725), .B(N5724), .S0(N3934));
MXI2XL addgen2_A_I1448 (.Y(N3943), .A(N5694), .B(N5693), .S0(N1103));
MXI2XL addgen2_A_I1449 (.Y(N1110), .A(N5725), .B(N5724), .S0(N3943));
MXI2XL addgen2_A_I1450 (.Y(N3952), .A(N5695), .B(N5694), .S0(N1103));
MXI2XL addgen2_A_I1451 (.Y(N1111), .A(N5725), .B(N5724), .S0(N3952));
MXI2XL addgen2_A_I1452 (.Y(N3961), .A(N5696), .B(N5695), .S0(N1103));
MXI2XL addgen2_A_I1453 (.Y(N1112), .A(N5725), .B(N5724), .S0(N3961));
MXI2XL addgen2_A_I1454 (.Y(N3970), .A(N5697), .B(N5696), .S0(N1103));
MXI2XL addgen2_A_I1455 (.Y(N1113), .A(N5725), .B(N5724), .S0(N3970));
MXI2XL addgen2_A_I1456 (.Y(N3979), .A(N5698), .B(N5697), .S0(N1103));
MXI2XL addgen2_A_I1457 (.Y(N1114), .A(N5725), .B(N5724), .S0(N3979));
MXI2XL addgen2_A_I1458 (.Y(N3988), .A(N5699), .B(N5698), .S0(N1103));
MXI2XL addgen2_A_I1459 (.Y(N1115), .A(N5725), .B(N5724), .S0(N3988));
MXI2XL addgen2_A_I1460 (.Y(N3997), .A(N5700), .B(N5699), .S0(N1103));
MXI2XL addgen2_A_I1461 (.Y(N1116), .A(N5725), .B(N5724), .S0(N3997));
MXI2XL addgen2_A_I1462 (.Y(N4006), .A(N5701), .B(N5700), .S0(N1103));
MXI2XL addgen2_A_I1463 (.Y(N1117), .A(N5725), .B(N5724), .S0(N4006));
MXI2XL addgen2_A_I1464 (.Y(N4015), .A(N5702), .B(N5701), .S0(N1103));
MXI2XL addgen2_A_I1465 (.Y(N1118), .A(N5725), .B(N5724), .S0(N4015));
MXI2XL addgen2_A_I1466 (.Y(N4024), .A(N5703), .B(N5702), .S0(N1103));
MXI2XL addgen2_A_I1467 (.Y(N1119), .A(N5725), .B(N5724), .S0(N4024));
MXI2XL addgen2_A_I1468 (.Y(N4033), .A(N5704), .B(N5703), .S0(N1103));
MXI2XL addgen2_A_I1469 (.Y(N1120), .A(N5725), .B(N5724), .S0(N4033));
MXI2XL addgen2_A_I1470 (.Y(N4042), .A(N5705), .B(N5704), .S0(N1103));
MXI2XL addgen2_A_I1471 (.Y(N1121), .A(N5725), .B(N5724), .S0(N4042));
MXI2XL addgen2_A_I1472 (.Y(N4051), .A(N5706), .B(N5705), .S0(N1103));
MXI2XL addgen2_A_I1473 (.Y(N1122), .A(N5725), .B(N5724), .S0(N4051));
MXI2XL addgen2_A_I1474 (.Y(N4060), .A(N5707), .B(N5706), .S0(N1103));
MXI2XL addgen2_A_I1475 (.Y(N1123), .A(N5725), .B(N5724), .S0(N4060));
MXI2XL addgen2_A_I1476 (.Y(N4069), .A(N5708), .B(N5707), .S0(N1103));
MXI2XL addgen2_A_I1477 (.Y(N1124), .A(N5725), .B(N5724), .S0(N4069));
MXI2XL addgen2_A_I1478 (.Y(N4078), .A(N5709), .B(N5708), .S0(N1103));
MXI2XL addgen2_A_I1479 (.Y(N1125), .A(N5725), .B(N5724), .S0(N4078));
MXI2XL addgen2_A_I1480 (.Y(N4087), .A(N5710), .B(N5709), .S0(N1103));
MXI2XL addgen2_A_I1481 (.Y(N1126), .A(N5725), .B(N5724), .S0(N4087));
MXI2XL addgen2_A_I1482 (.Y(N4096), .A(N5711), .B(N5710), .S0(N1103));
MXI2XL addgen2_A_I1483 (.Y(N1127), .A(N5725), .B(N5724), .S0(N4096));
MXI2XL addgen2_A_I1484 (.Y(N4105), .A(N5712), .B(N5711), .S0(N1103));
MXI2XL addgen2_A_I1485 (.Y(N1128), .A(N5725), .B(N5724), .S0(N4105));
MXI2XL addgen2_A_I1486 (.Y(N4114), .A(N5713), .B(N5712), .S0(N1103));
MXI2XL addgen2_A_I1487 (.Y(N1129), .A(N5725), .B(N5724), .S0(N4114));
MXI2XL addgen2_A_I1488 (.Y(N4123), .A(N5714), .B(N5713), .S0(N1103));
MXI2XL addgen2_A_I1489 (.Y(N1130), .A(N5725), .B(N5724), .S0(N4123));
NOR2BX1 addgen2_A_I1490 (.Y(N4132), .AN(N1103), .B(N5714));
MXI2XL addgen2_A_I1491 (.Y(N1131), .A(N5725), .B(N5724), .S0(N4132));
XNOR2X1 enc2_A_I1492 (.Y(N1135), .A(inst_cellmath__203_0_in0[5]), .B(inst_cellmath__203_0_in0[4]));
NOR2XL enc2_A_I1494 (.Y(N4143), .A(inst_cellmath__203_0_in0[5]), .B(inst_cellmath__203_0_in0[4]));
OAI2BB1X1 enc2_A_I1833 (.Y(N1134), .A0N(inst_cellmath__203_0_in0[5]), .A1N(inst_cellmath__203_0_in0[4]), .B0(inst_cellmath__203_0_in0[6]));
INVXL inst_cellmath__203_0_I1930 (.Y(N5726), .A(N1134));
OR2XL inst_cellmath__203_0_I1977 (.Y(N5729), .A(N4143), .B(inst_cellmath__203_0_in0[6]));
INVXL inst_cellmath__203_0_I1934 (.Y(N5730), .A(N5726));
NOR2XL addgen2_A_I1497 (.Y(N4154), .A(N5693), .B(N1135));
MXI2XL addgen2_A_I1498 (.Y(N1141), .A(N5730), .B(N5729), .S0(N4154));
MXI2XL addgen2_A_I1499 (.Y(N4163), .A(N5694), .B(N5693), .S0(N1135));
MXI2XL addgen2_A_I1500 (.Y(N1142), .A(N5730), .B(N5729), .S0(N4163));
MXI2XL addgen2_A_I1501 (.Y(N4172), .A(N5695), .B(N5694), .S0(N1135));
MXI2XL addgen2_A_I1502 (.Y(N1143), .A(N5730), .B(N5729), .S0(N4172));
MXI2XL addgen2_A_I1503 (.Y(N4181), .A(N5696), .B(N5695), .S0(N1135));
MXI2XL addgen2_A_I1504 (.Y(N1144), .A(N5730), .B(N5729), .S0(N4181));
MXI2XL addgen2_A_I1505 (.Y(N4190), .A(N5697), .B(N5696), .S0(N1135));
MXI2XL addgen2_A_I1506 (.Y(N1145), .A(N5730), .B(N5729), .S0(N4190));
MXI2XL addgen2_A_I1507 (.Y(N4199), .A(N5698), .B(N5697), .S0(N1135));
MXI2XL addgen2_A_I1508 (.Y(N1146), .A(N5730), .B(N5729), .S0(N4199));
MXI2XL addgen2_A_I1509 (.Y(N4208), .A(N5699), .B(N5698), .S0(N1135));
MXI2XL addgen2_A_I1510 (.Y(N1147), .A(N5730), .B(N5729), .S0(N4208));
MXI2XL addgen2_A_I1511 (.Y(N4217), .A(N5700), .B(N5699), .S0(N1135));
MXI2XL addgen2_A_I1512 (.Y(N1148), .A(N5730), .B(N5729), .S0(N4217));
MXI2XL addgen2_A_I1513 (.Y(N4226), .A(N5701), .B(N5700), .S0(N1135));
MXI2XL addgen2_A_I1514 (.Y(N1149), .A(N5730), .B(N5729), .S0(N4226));
MXI2XL addgen2_A_I1515 (.Y(N4235), .A(N5702), .B(N5701), .S0(N1135));
MXI2XL addgen2_A_I1516 (.Y(N1150), .A(N5730), .B(N5729), .S0(N4235));
MXI2XL addgen2_A_I1517 (.Y(N4244), .A(N5703), .B(N5702), .S0(N1135));
MXI2XL addgen2_A_I1518 (.Y(N1151), .A(N5730), .B(N5729), .S0(N4244));
MXI2XL addgen2_A_I1519 (.Y(N4253), .A(N5704), .B(N5703), .S0(N1135));
MXI2XL addgen2_A_I1520 (.Y(N1152), .A(N5730), .B(N5729), .S0(N4253));
MXI2XL addgen2_A_I1521 (.Y(N4262), .A(N5705), .B(N5704), .S0(N1135));
MXI2XL addgen2_A_I1522 (.Y(N1153), .A(N5730), .B(N5729), .S0(N4262));
MXI2XL addgen2_A_I1523 (.Y(N4271), .A(N5706), .B(N5705), .S0(N1135));
MXI2XL addgen2_A_I1524 (.Y(N1154), .A(N5730), .B(N5729), .S0(N4271));
MXI2XL addgen2_A_I1525 (.Y(N4280), .A(N5707), .B(N5706), .S0(N1135));
MXI2XL addgen2_A_I1526 (.Y(N1155), .A(N5730), .B(N5729), .S0(N4280));
MXI2XL addgen2_A_I1527 (.Y(N4289), .A(N5708), .B(N5707), .S0(N1135));
MXI2XL addgen2_A_I1528 (.Y(N1156), .A(N5730), .B(N5729), .S0(N4289));
MXI2XL addgen2_A_I1529 (.Y(N4298), .A(N5709), .B(N5708), .S0(N1135));
MXI2XL addgen2_A_I1530 (.Y(N1157), .A(N5730), .B(N5729), .S0(N4298));
MXI2XL addgen2_A_I1531 (.Y(N4307), .A(N5710), .B(N5709), .S0(N1135));
MXI2XL addgen2_A_I1532 (.Y(N1158), .A(N5730), .B(N5729), .S0(N4307));
MXI2XL addgen2_A_I1533 (.Y(N4316), .A(N5711), .B(N5710), .S0(N1135));
MXI2XL addgen2_A_I1534 (.Y(N1159), .A(N5730), .B(N5729), .S0(N4316));
MXI2XL addgen2_A_I1535 (.Y(N4325), .A(N5712), .B(N5711), .S0(N1135));
MXI2XL addgen2_A_I1536 (.Y(N1160), .A(N5730), .B(N5729), .S0(N4325));
MXI2XL addgen2_A_I1537 (.Y(N4334), .A(N5713), .B(N5712), .S0(N1135));
MXI2XL addgen2_A_I1538 (.Y(N1161), .A(N5730), .B(N5729), .S0(N4334));
MXI2XL addgen2_A_I1539 (.Y(N4343), .A(N5714), .B(N5713), .S0(N1135));
MXI2XL addgen2_A_I1540 (.Y(N1162), .A(N5730), .B(N5729), .S0(N4343));
NOR2BX1 addgen2_A_I1541 (.Y(N4352), .AN(N1135), .B(N5714));
MXI2XL addgen2_A_I1542 (.Y(N1163), .A(N5730), .B(N5729), .S0(N4352));
XNOR2X1 enc2_A_I1543 (.Y(N1167), .A(inst_cellmath__203_0_in0[7]), .B(inst_cellmath__203_0_in0[6]));
NOR2XL enc2_A_I1545 (.Y(N4363), .A(inst_cellmath__203_0_in0[7]), .B(inst_cellmath__203_0_in0[6]));
OAI2BB1X1 enc2_A_I1834 (.Y(N1166), .A0N(inst_cellmath__203_0_in0[7]), .A1N(inst_cellmath__203_0_in0[6]), .B0(inst_cellmath__203_0_in0[8]));
INVXL inst_cellmath__203_0_I1935 (.Y(N5731), .A(N1166));
OR2XL inst_cellmath__203_0_I1978 (.Y(N5734), .A(N4363), .B(inst_cellmath__203_0_in0[8]));
INVXL inst_cellmath__203_0_I1939 (.Y(N5735), .A(N5731));
NOR2XL addgen2_A_I1548 (.Y(N4374), .A(N5693), .B(N1167));
MXI2XL addgen2_A_I1549 (.Y(N1173), .A(N5735), .B(N5734), .S0(N4374));
MXI2XL addgen2_A_I1550 (.Y(N4383), .A(N5694), .B(N5693), .S0(N1167));
MXI2XL addgen2_A_I1551 (.Y(N1174), .A(N5735), .B(N5734), .S0(N4383));
MXI2XL addgen2_A_I1552 (.Y(N4392), .A(N5695), .B(N5694), .S0(N1167));
MXI2XL addgen2_A_I1553 (.Y(N1175), .A(N5735), .B(N5734), .S0(N4392));
MXI2XL addgen2_A_I1554 (.Y(N4401), .A(N5696), .B(N5695), .S0(N1167));
MXI2XL addgen2_A_I1555 (.Y(N1176), .A(N5735), .B(N5734), .S0(N4401));
MXI2XL addgen2_A_I1556 (.Y(N4410), .A(N5697), .B(N5696), .S0(N1167));
MXI2XL addgen2_A_I1557 (.Y(N1177), .A(N5735), .B(N5734), .S0(N4410));
MXI2XL addgen2_A_I1558 (.Y(N4419), .A(N5698), .B(N5697), .S0(N1167));
MXI2XL addgen2_A_I1559 (.Y(N1178), .A(N5735), .B(N5734), .S0(N4419));
MXI2XL addgen2_A_I1560 (.Y(N4428), .A(N5699), .B(N5698), .S0(N1167));
MXI2XL addgen2_A_I1561 (.Y(N1179), .A(N5735), .B(N5734), .S0(N4428));
MXI2XL addgen2_A_I1562 (.Y(N4437), .A(N5700), .B(N5699), .S0(N1167));
MXI2XL addgen2_A_I1563 (.Y(N1180), .A(N5735), .B(N5734), .S0(N4437));
MXI2XL addgen2_A_I1564 (.Y(N4446), .A(N5701), .B(N5700), .S0(N1167));
MXI2XL addgen2_A_I1565 (.Y(N1181), .A(N5735), .B(N5734), .S0(N4446));
MXI2XL addgen2_A_I1566 (.Y(N4455), .A(N5702), .B(N5701), .S0(N1167));
MXI2XL addgen2_A_I1567 (.Y(N1182), .A(N5735), .B(N5734), .S0(N4455));
MXI2XL addgen2_A_I1568 (.Y(N4464), .A(N5703), .B(N5702), .S0(N1167));
MXI2XL addgen2_A_I1569 (.Y(N1183), .A(N5735), .B(N5734), .S0(N4464));
MXI2XL addgen2_A_I1570 (.Y(N4473), .A(N5704), .B(N5703), .S0(N1167));
MXI2XL addgen2_A_I1571 (.Y(N1184), .A(N5735), .B(N5734), .S0(N4473));
MXI2XL addgen2_A_I1572 (.Y(N4482), .A(N5705), .B(N5704), .S0(N1167));
MXI2XL addgen2_A_I1573 (.Y(N1185), .A(N5735), .B(N5734), .S0(N4482));
MXI2XL addgen2_A_I1574 (.Y(N4491), .A(N5706), .B(N5705), .S0(N1167));
MXI2XL addgen2_A_I1575 (.Y(N1186), .A(N5735), .B(N5734), .S0(N4491));
MXI2XL addgen2_A_I1576 (.Y(N4500), .A(N5707), .B(N5706), .S0(N1167));
MXI2XL addgen2_A_I1577 (.Y(N1187), .A(N5735), .B(N5734), .S0(N4500));
MXI2XL addgen2_A_I1578 (.Y(N4509), .A(N5708), .B(N5707), .S0(N1167));
MXI2XL addgen2_A_I1579 (.Y(N1188), .A(N5735), .B(N5734), .S0(N4509));
MXI2XL addgen2_A_I1580 (.Y(N4518), .A(N5709), .B(N5708), .S0(N1167));
MXI2XL addgen2_A_I1581 (.Y(N1189), .A(N5735), .B(N5734), .S0(N4518));
MXI2XL addgen2_A_I1582 (.Y(N4527), .A(N5710), .B(N5709), .S0(N1167));
MXI2XL addgen2_A_I1583 (.Y(N1190), .A(N5735), .B(N5734), .S0(N4527));
MXI2XL addgen2_A_I1584 (.Y(N4536), .A(N5711), .B(N5710), .S0(N1167));
MXI2XL addgen2_A_I1585 (.Y(N1191), .A(N5735), .B(N5734), .S0(N4536));
MXI2XL addgen2_A_I1586 (.Y(N4545), .A(N5712), .B(N5711), .S0(N1167));
MXI2XL addgen2_A_I1587 (.Y(N1192), .A(N5735), .B(N5734), .S0(N4545));
MXI2XL addgen2_A_I1588 (.Y(N4554), .A(N5713), .B(N5712), .S0(N1167));
MXI2XL addgen2_A_I1589 (.Y(N1193), .A(N5735), .B(N5734), .S0(N4554));
MXI2XL addgen2_A_I1590 (.Y(N4563), .A(N5714), .B(N5713), .S0(N1167));
MXI2XL addgen2_A_I1591 (.Y(N1194), .A(N5735), .B(N5734), .S0(N4563));
NOR2BX1 addgen2_A_I1592 (.Y(N4572), .AN(N1167), .B(N5714));
MXI2XL addgen2_A_I1593 (.Y(N1195), .A(N5735), .B(N5734), .S0(N4572));
XNOR2X1 enc2_A_I1594 (.Y(N1199), .A(inst_cellmath__203_0_in0[9]), .B(inst_cellmath__203_0_in0[8]));
NOR2XL enc2_A_I1596 (.Y(N4583), .A(inst_cellmath__203_0_in0[9]), .B(inst_cellmath__203_0_in0[8]));
OAI2BB1X1 enc2_A_I1835 (.Y(N1198), .A0N(inst_cellmath__203_0_in0[9]), .A1N(inst_cellmath__203_0_in0[8]), .B0(inst_cellmath__203_0_in0[10]));
INVXL inst_cellmath__203_0_I1940 (.Y(N5736), .A(N1198));
OR2XL inst_cellmath__203_0_I1979 (.Y(N5739), .A(N4583), .B(inst_cellmath__203_0_in0[10]));
INVXL inst_cellmath__203_0_I1944 (.Y(N5740), .A(N5736));
NOR2XL addgen2_A_I1599 (.Y(N4594), .A(N5693), .B(N1199));
MXI2XL addgen2_A_I1600 (.Y(N1205), .A(N5740), .B(N5739), .S0(N4594));
MXI2XL addgen2_A_I1601 (.Y(N4603), .A(N5694), .B(N5693), .S0(N1199));
MXI2XL addgen2_A_I1602 (.Y(N1206), .A(N5740), .B(N5739), .S0(N4603));
MXI2XL addgen2_A_I1603 (.Y(N4612), .A(N5695), .B(N5694), .S0(N1199));
MXI2XL addgen2_A_I1604 (.Y(N1207), .A(N5740), .B(N5739), .S0(N4612));
MXI2XL addgen2_A_I1605 (.Y(N4621), .A(N5696), .B(N5695), .S0(N1199));
MXI2XL addgen2_A_I1606 (.Y(N1208), .A(N5740), .B(N5739), .S0(N4621));
MXI2XL addgen2_A_I1607 (.Y(N4630), .A(N5697), .B(N5696), .S0(N1199));
MXI2XL addgen2_A_I1608 (.Y(N1209), .A(N5740), .B(N5739), .S0(N4630));
MXI2XL addgen2_A_I1609 (.Y(N4639), .A(N5698), .B(N5697), .S0(N1199));
MXI2XL addgen2_A_I1610 (.Y(N1210), .A(N5740), .B(N5739), .S0(N4639));
MXI2XL addgen2_A_I1611 (.Y(N4648), .A(N5699), .B(N5698), .S0(N1199));
MXI2XL addgen2_A_I1612 (.Y(N1211), .A(N5740), .B(N5739), .S0(N4648));
MXI2XL addgen2_A_I1613 (.Y(N4657), .A(N5700), .B(N5699), .S0(N1199));
MXI2XL addgen2_A_I1614 (.Y(N1212), .A(N5740), .B(N5739), .S0(N4657));
MXI2XL addgen2_A_I1615 (.Y(N4666), .A(N5701), .B(N5700), .S0(N1199));
MXI2XL addgen2_A_I1616 (.Y(N1213), .A(N5740), .B(N5739), .S0(N4666));
MXI2XL addgen2_A_I1617 (.Y(N4675), .A(N5702), .B(N5701), .S0(N1199));
MXI2XL addgen2_A_I1618 (.Y(N1214), .A(N5740), .B(N5739), .S0(N4675));
MXI2XL addgen2_A_I1619 (.Y(N4684), .A(N5703), .B(N5702), .S0(N1199));
MXI2XL addgen2_A_I1620 (.Y(N1215), .A(N5740), .B(N5739), .S0(N4684));
MXI2XL addgen2_A_I1621 (.Y(N4693), .A(N5704), .B(N5703), .S0(N1199));
MXI2XL addgen2_A_I1622 (.Y(N1216), .A(N5740), .B(N5739), .S0(N4693));
MXI2XL addgen2_A_I1623 (.Y(N4702), .A(N5705), .B(N5704), .S0(N1199));
MXI2XL addgen2_A_I1624 (.Y(N1217), .A(N5740), .B(N5739), .S0(N4702));
MXI2XL addgen2_A_I1625 (.Y(N4711), .A(N5706), .B(N5705), .S0(N1199));
MXI2XL addgen2_A_I1626 (.Y(N1218), .A(N5740), .B(N5739), .S0(N4711));
MXI2XL addgen2_A_I1627 (.Y(N4720), .A(N5707), .B(N5706), .S0(N1199));
MXI2XL addgen2_A_I1628 (.Y(N1219), .A(N5740), .B(N5739), .S0(N4720));
MXI2XL addgen2_A_I1629 (.Y(N4729), .A(N5708), .B(N5707), .S0(N1199));
MXI2XL addgen2_A_I1630 (.Y(N1220), .A(N5740), .B(N5739), .S0(N4729));
MXI2XL addgen2_A_I1631 (.Y(N4738), .A(N5709), .B(N5708), .S0(N1199));
MXI2XL addgen2_A_I1632 (.Y(N1221), .A(N5740), .B(N5739), .S0(N4738));
MXI2XL addgen2_A_I1633 (.Y(N4747), .A(N5710), .B(N5709), .S0(N1199));
MXI2XL addgen2_A_I1634 (.Y(N1222), .A(N5740), .B(N5739), .S0(N4747));
MXI2XL addgen2_A_I1635 (.Y(N4756), .A(N5711), .B(N5710), .S0(N1199));
MXI2XL addgen2_A_I1636 (.Y(N1223), .A(N5740), .B(N5739), .S0(N4756));
MXI2XL addgen2_A_I1637 (.Y(N4765), .A(N5712), .B(N5711), .S0(N1199));
MXI2XL addgen2_A_I1638 (.Y(N1224), .A(N5740), .B(N5739), .S0(N4765));
MXI2XL addgen2_A_I1639 (.Y(N4774), .A(N5713), .B(N5712), .S0(N1199));
MXI2XL addgen2_A_I1640 (.Y(N1225), .A(N5740), .B(N5739), .S0(N4774));
MXI2XL addgen2_A_I1641 (.Y(N4783), .A(N5714), .B(N5713), .S0(N1199));
MXI2XL addgen2_A_I1642 (.Y(N1226), .A(N5740), .B(N5739), .S0(N4783));
NOR2BX1 addgen2_A_I1643 (.Y(N4792), .AN(N1199), .B(N5714));
MXI2XL addgen2_A_I1644 (.Y(N1227), .A(N5740), .B(N5739), .S0(N4792));
XNOR2X1 enc2_A_I1645 (.Y(N1231), .A(inst_cellmath__203_0_in0[11]), .B(inst_cellmath__203_0_in0[10]));
NOR2XL enc2_A_I1647 (.Y(N4803), .A(inst_cellmath__203_0_in0[11]), .B(inst_cellmath__203_0_in0[10]));
OAI2BB1X1 enc2_A_I1836 (.Y(N1230), .A0N(inst_cellmath__203_0_in0[11]), .A1N(inst_cellmath__203_0_in0[10]), .B0(inst_cellmath__203_0_in0[12]));
INVXL inst_cellmath__203_0_I1945 (.Y(N5741), .A(N1230));
OR2XL inst_cellmath__203_0_I1980 (.Y(N5744), .A(N4803), .B(inst_cellmath__203_0_in0[12]));
INVXL inst_cellmath__203_0_I1949 (.Y(N5745), .A(N5741));
NOR2XL addgen2_A_I1650 (.Y(N4814), .A(N5693), .B(N1231));
MXI2XL addgen2_A_I1651 (.Y(N1237), .A(N5745), .B(N5744), .S0(N4814));
MXI2XL addgen2_A_I1652 (.Y(N4823), .A(N5694), .B(N5693), .S0(N1231));
MXI2XL addgen2_A_I1653 (.Y(N1238), .A(N5745), .B(N5744), .S0(N4823));
MXI2XL addgen2_A_I1654 (.Y(N4832), .A(N5695), .B(N5694), .S0(N1231));
MXI2XL addgen2_A_I1655 (.Y(N1239), .A(N5745), .B(N5744), .S0(N4832));
MXI2XL addgen2_A_I1656 (.Y(N4841), .A(N5696), .B(N5695), .S0(N1231));
MXI2XL addgen2_A_I1657 (.Y(N1240), .A(N5745), .B(N5744), .S0(N4841));
MXI2XL addgen2_A_I1658 (.Y(N4850), .A(N5697), .B(N5696), .S0(N1231));
MXI2XL addgen2_A_I1659 (.Y(N1241), .A(N5745), .B(N5744), .S0(N4850));
MXI2XL addgen2_A_I1660 (.Y(N4859), .A(N5698), .B(N5697), .S0(N1231));
MXI2XL addgen2_A_I1661 (.Y(N1242), .A(N5745), .B(N5744), .S0(N4859));
MXI2XL addgen2_A_I1662 (.Y(N4868), .A(N5699), .B(N5698), .S0(N1231));
MXI2XL addgen2_A_I1663 (.Y(N1243), .A(N5745), .B(N5744), .S0(N4868));
MXI2XL addgen2_A_I1664 (.Y(N4877), .A(N5700), .B(N5699), .S0(N1231));
MXI2XL addgen2_A_I1665 (.Y(N1244), .A(N5745), .B(N5744), .S0(N4877));
MXI2XL addgen2_A_I1666 (.Y(N4886), .A(N5701), .B(N5700), .S0(N1231));
MXI2XL addgen2_A_I1667 (.Y(N1245), .A(N5745), .B(N5744), .S0(N4886));
MXI2XL addgen2_A_I1668 (.Y(N4895), .A(N5702), .B(N5701), .S0(N1231));
MXI2XL addgen2_A_I1669 (.Y(N1246), .A(N5745), .B(N5744), .S0(N4895));
MXI2XL addgen2_A_I1670 (.Y(N4904), .A(N5703), .B(N5702), .S0(N1231));
MXI2XL addgen2_A_I1671 (.Y(N1247), .A(N5745), .B(N5744), .S0(N4904));
MXI2XL addgen2_A_I1672 (.Y(N4913), .A(N5704), .B(N5703), .S0(N1231));
MXI2XL addgen2_A_I1673 (.Y(N1248), .A(N5745), .B(N5744), .S0(N4913));
MXI2XL addgen2_A_I1674 (.Y(N4922), .A(N5705), .B(N5704), .S0(N1231));
MXI2XL addgen2_A_I1675 (.Y(N1249), .A(N5745), .B(N5744), .S0(N4922));
MXI2XL addgen2_A_I1676 (.Y(N4931), .A(N5706), .B(N5705), .S0(N1231));
MXI2XL addgen2_A_I1677 (.Y(N1250), .A(N5745), .B(N5744), .S0(N4931));
MXI2XL addgen2_A_I1678 (.Y(N4940), .A(N5707), .B(N5706), .S0(N1231));
MXI2XL addgen2_A_I1679 (.Y(N1251), .A(N5745), .B(N5744), .S0(N4940));
MXI2XL addgen2_A_I1680 (.Y(N4949), .A(N5708), .B(N5707), .S0(N1231));
MXI2XL addgen2_A_I1681 (.Y(N1252), .A(N5745), .B(N5744), .S0(N4949));
MXI2XL addgen2_A_I1682 (.Y(N4958), .A(N5709), .B(N5708), .S0(N1231));
MXI2XL addgen2_A_I1683 (.Y(N1253), .A(N5745), .B(N5744), .S0(N4958));
MXI2XL addgen2_A_I1684 (.Y(N4967), .A(N5710), .B(N5709), .S0(N1231));
MXI2XL addgen2_A_I1685 (.Y(N1254), .A(N5745), .B(N5744), .S0(N4967));
MXI2XL addgen2_A_I1686 (.Y(N4976), .A(N5711), .B(N5710), .S0(N1231));
MXI2XL addgen2_A_I1687 (.Y(N1255), .A(N5745), .B(N5744), .S0(N4976));
MXI2XL addgen2_A_I1688 (.Y(N4985), .A(N5712), .B(N5711), .S0(N1231));
MXI2XL addgen2_A_I1689 (.Y(N1256), .A(N5745), .B(N5744), .S0(N4985));
MXI2XL addgen2_A_I1690 (.Y(N4994), .A(N5713), .B(N5712), .S0(N1231));
MXI2XL addgen2_A_I1691 (.Y(N1257), .A(N5745), .B(N5744), .S0(N4994));
MXI2XL addgen2_A_I1692 (.Y(N5003), .A(N5714), .B(N5713), .S0(N1231));
MXI2XL addgen2_A_I1693 (.Y(N1258), .A(N5745), .B(N5744), .S0(N5003));
NOR2BX1 addgen2_A_I1694 (.Y(N5012), .AN(N1231), .B(N5714));
MXI2XL addgen2_A_I1695 (.Y(N1259), .A(N5745), .B(N5744), .S0(N5012));
XNOR2X1 enc2_A_I1696 (.Y(N1263), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
NOR2XL enc2_A_I1698 (.Y(N5023), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
OAI2BB1X1 enc2_A_I1837 (.Y(N1262), .A0N(inst_cellmath__203_0_in0[13]), .A1N(inst_cellmath__203_0_in0[12]), .B0(inst_cellmath__203_0_in0[14]));
INVXL inst_cellmath__203_0_I1950 (.Y(N5746), .A(N1262));
OR2XL inst_cellmath__203_0_I1981 (.Y(N5749), .A(N5023), .B(inst_cellmath__203_0_in0[14]));
INVXL inst_cellmath__203_0_I1954 (.Y(N5750), .A(N5746));
NOR2XL addgen2_A_I1701 (.Y(N5034), .A(N5693), .B(N1263));
MXI2XL addgen2_A_I1702 (.Y(N1269), .A(N5750), .B(N5749), .S0(N5034));
MXI2XL addgen2_A_I1703 (.Y(N5043), .A(N5694), .B(N5693), .S0(N1263));
MXI2XL addgen2_A_I1704 (.Y(N1270), .A(N5750), .B(N5749), .S0(N5043));
MXI2XL addgen2_A_I1705 (.Y(N5052), .A(N5695), .B(N5694), .S0(N1263));
MXI2XL addgen2_A_I1706 (.Y(N1271), .A(N5750), .B(N5749), .S0(N5052));
MXI2XL addgen2_A_I1707 (.Y(N5061), .A(N5696), .B(N5695), .S0(N1263));
MXI2XL addgen2_A_I1708 (.Y(N1272), .A(N5750), .B(N5749), .S0(N5061));
MXI2XL addgen2_A_I1709 (.Y(N5070), .A(N5697), .B(N5696), .S0(N1263));
MXI2XL addgen2_A_I1710 (.Y(N1273), .A(N5750), .B(N5749), .S0(N5070));
MXI2XL addgen2_A_I1711 (.Y(N5079), .A(N5698), .B(N5697), .S0(N1263));
MXI2XL addgen2_A_I1712 (.Y(N1274), .A(N5750), .B(N5749), .S0(N5079));
MXI2XL addgen2_A_I1713 (.Y(N5088), .A(N5699), .B(N5698), .S0(N1263));
MXI2XL addgen2_A_I1714 (.Y(N1275), .A(N5750), .B(N5749), .S0(N5088));
MXI2XL addgen2_A_I1715 (.Y(N5097), .A(N5700), .B(N5699), .S0(N1263));
MXI2XL addgen2_A_I1716 (.Y(N1276), .A(N5750), .B(N5749), .S0(N5097));
MXI2XL addgen2_A_I1717 (.Y(N5106), .A(N5701), .B(N5700), .S0(N1263));
MXI2XL addgen2_A_I1718 (.Y(N1277), .A(N5750), .B(N5749), .S0(N5106));
MXI2XL addgen2_A_I1719 (.Y(N5115), .A(N5702), .B(N5701), .S0(N1263));
MXI2XL addgen2_A_I1720 (.Y(N1278), .A(N5750), .B(N5749), .S0(N5115));
MXI2XL addgen2_A_I1721 (.Y(N5124), .A(N5703), .B(N5702), .S0(N1263));
MXI2XL addgen2_A_I1722 (.Y(N1279), .A(N5750), .B(N5749), .S0(N5124));
MXI2XL addgen2_A_I1723 (.Y(N5133), .A(N5704), .B(N5703), .S0(N1263));
MXI2XL addgen2_A_I1724 (.Y(N1280), .A(N5750), .B(N5749), .S0(N5133));
MXI2XL addgen2_A_I1725 (.Y(N5142), .A(N5705), .B(N5704), .S0(N1263));
MXI2XL addgen2_A_I1726 (.Y(N1281), .A(N5750), .B(N5749), .S0(N5142));
MXI2XL addgen2_A_I1727 (.Y(N5151), .A(N5706), .B(N5705), .S0(N1263));
MXI2XL addgen2_A_I1728 (.Y(N1282), .A(N5750), .B(N5749), .S0(N5151));
MXI2XL addgen2_A_I1729 (.Y(N5160), .A(N5707), .B(N5706), .S0(N1263));
MXI2XL addgen2_A_I1730 (.Y(N1283), .A(N5750), .B(N5749), .S0(N5160));
MXI2XL addgen2_A_I1731 (.Y(N5169), .A(N5708), .B(N5707), .S0(N1263));
MXI2XL addgen2_A_I1732 (.Y(N1284), .A(N5750), .B(N5749), .S0(N5169));
MXI2XL addgen2_A_I1733 (.Y(N5178), .A(N5709), .B(N5708), .S0(N1263));
MXI2XL addgen2_A_I1734 (.Y(N1285), .A(N5750), .B(N5749), .S0(N5178));
MXI2XL addgen2_A_I1735 (.Y(N5187), .A(N5710), .B(N5709), .S0(N1263));
MXI2XL addgen2_A_I1736 (.Y(N1286), .A(N5750), .B(N5749), .S0(N5187));
MXI2XL addgen2_A_I1737 (.Y(N5196), .A(N5711), .B(N5710), .S0(N1263));
MXI2XL addgen2_A_I1738 (.Y(N1287), .A(N5750), .B(N5749), .S0(N5196));
MXI2XL addgen2_A_I1739 (.Y(N5205), .A(N5712), .B(N5711), .S0(N1263));
MXI2XL addgen2_A_I1740 (.Y(N1288), .A(N5750), .B(N5749), .S0(N5205));
MXI2XL addgen2_A_I1741 (.Y(N5214), .A(N5713), .B(N5712), .S0(N1263));
MXI2XL addgen2_A_I1742 (.Y(N1289), .A(N5750), .B(N5749), .S0(N5214));
MXI2XL addgen2_A_I1743 (.Y(N5223), .A(N5714), .B(N5713), .S0(N1263));
MXI2XL addgen2_A_I1744 (.Y(N1290), .A(N5750), .B(N5749), .S0(N5223));
NOR2BX1 addgen2_A_I1745 (.Y(N5232), .AN(N1263), .B(N5714));
MXI2XL addgen2_A_I1746 (.Y(N2112), .A(N5750), .B(N5749), .S0(N5232));
XNOR2X1 enc2_A_I1747 (.Y(N1295), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
NOR2XL enc2_A_I1749 (.Y(N5243), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
OAI2BB1X1 enc2_A_I1838 (.Y(N1294), .A0N(inst_cellmath__203_0_in0[15]), .A1N(inst_cellmath__203_0_in0[14]), .B0(inst_cellmath__203_0_in4[0]));
INVXL inst_cellmath__203_0_I1955 (.Y(N5751), .A(N1294));
OR2XL inst_cellmath__203_0_I1982 (.Y(N5754), .A(N5243), .B(inst_cellmath__203_0_in4[0]));
INVXL inst_cellmath__203_0_I1959 (.Y(inst_cellmath__203_0_out1[42]), .A(N5751));
NOR2XL addgen2_A_I1752 (.Y(N5254), .A(N5693), .B(N1295));
MXI2XL addgen2_A_I1753 (.Y(N1301), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5254));
MXI2XL addgen2_A_I1754 (.Y(N5263), .A(N5694), .B(N5693), .S0(N1295));
MXI2XL addgen2_A_I1755 (.Y(N1302), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5263));
MXI2XL addgen2_A_I1756 (.Y(N5272), .A(N5695), .B(N5694), .S0(N1295));
MXI2XL addgen2_A_I1757 (.Y(N1303), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5272));
MXI2XL addgen2_A_I1758 (.Y(N5281), .A(N5696), .B(N5695), .S0(N1295));
MXI2XL addgen2_A_I1759 (.Y(N1304), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5281));
MXI2XL addgen2_A_I1760 (.Y(N5290), .A(N5697), .B(N5696), .S0(N1295));
MXI2XL addgen2_A_I1761 (.Y(N1305), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5290));
MXI2XL addgen2_A_I1762 (.Y(N5299), .A(N5698), .B(N5697), .S0(N1295));
MXI2XL addgen2_A_I1763 (.Y(N1306), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5299));
MXI2XL addgen2_A_I1764 (.Y(N5308), .A(N5699), .B(N5698), .S0(N1295));
MXI2XL addgen2_A_I1765 (.Y(N1307), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5308));
MXI2XL addgen2_A_I1766 (.Y(N5317), .A(N5700), .B(N5699), .S0(N1295));
MXI2XL addgen2_A_I1767 (.Y(N1308), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5317));
MXI2XL addgen2_A_I1768 (.Y(N5326), .A(N5701), .B(N5700), .S0(N1295));
MXI2XL addgen2_A_I1769 (.Y(N1309), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5326));
MXI2XL addgen2_A_I1770 (.Y(N5335), .A(N5702), .B(N5701), .S0(N1295));
MXI2XL addgen2_A_I1771 (.Y(N1310), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5335));
MXI2XL addgen2_A_I1772 (.Y(N5344), .A(N5703), .B(N5702), .S0(N1295));
MXI2XL addgen2_A_I1773 (.Y(N1311), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5344));
MXI2XL addgen2_A_I1774 (.Y(N5353), .A(N5704), .B(N5703), .S0(N1295));
MXI2XL addgen2_A_I1775 (.Y(N1312), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5353));
MXI2XL addgen2_A_I1776 (.Y(N5362), .A(N5705), .B(N5704), .S0(N1295));
MXI2XL addgen2_A_I1777 (.Y(N1313), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5362));
MXI2XL addgen2_A_I1778 (.Y(N5371), .A(N5706), .B(N5705), .S0(N1295));
MXI2XL addgen2_A_I1779 (.Y(N1314), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5371));
MXI2XL addgen2_A_I1780 (.Y(N5380), .A(N5707), .B(N5706), .S0(N1295));
MXI2XL addgen2_A_I1781 (.Y(N1315), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5380));
MXI2XL addgen2_A_I1782 (.Y(N5389), .A(N5708), .B(N5707), .S0(N1295));
MXI2XL addgen2_A_I1783 (.Y(N1316), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5389));
MXI2XL addgen2_A_I1784 (.Y(N5398), .A(N5709), .B(N5708), .S0(N1295));
MXI2XL addgen2_A_I1785 (.Y(N1317), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5398));
MXI2XL addgen2_A_I1786 (.Y(N5407), .A(N5710), .B(N5709), .S0(N1295));
MXI2XL addgen2_A_I1787 (.Y(N1318), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5407));
MXI2XL addgen2_A_I1788 (.Y(N5416), .A(N5711), .B(N5710), .S0(N1295));
MXI2XL addgen2_A_I1789 (.Y(N1319), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5416));
MXI2XL addgen2_A_I1790 (.Y(N5425), .A(N5712), .B(N5711), .S0(N1295));
MXI2XL addgen2_A_I1791 (.Y(N1320), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5425));
MXI2XL addgen2_A_I1792 (.Y(N5434), .A(N5713), .B(N5712), .S0(N1295));
MXI2XL addgen2_A_I1793 (.Y(N1321), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5434));
MXI2XL addgen2_A_I1794 (.Y(N5443), .A(N5714), .B(N5713), .S0(N1295));
MXI2XL addgen2_A_I1795 (.Y(N1322), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5443));
NOR2BX1 addgen2_A_I1796 (.Y(N5452), .AN(N1295), .B(N5714));
MXI2XL addgen2_A_I1797 (.Y(inst_cellmath__203_0_out0[42]), .A(inst_cellmath__203_0_out1[42]), .B(N5754), .S0(N5452));
ADDHX1 inst_cellmath__203_0_I684 (.CO(inst_cellmath__203_0_out1[2]), .S(inst_cellmath__203_0_out0[1]), .A(N518), .B(inst_cellmath__203_0_in1[19]));
ADDHX1 inst_cellmath__203_0_I685 (.CO(inst_cellmath__203_0_out1[3]), .S(inst_cellmath__203_0_out0[2]), .A(N520), .B(N566));
ADDHX1 inst_cellmath__203_0_I686 (.CO(N1380), .S(N1379), .A(N522), .B(N5661));
ADDFX1 inst_cellmath__203_0_I687 (.CO(inst_cellmath__203_0_out1[4]), .S(inst_cellmath__203_0_out0[3]), .A(N595), .B(N567), .CI(N1379));
ADDFX1 inst_cellmath__203_0_I688 (.CO(N1384), .S(N1383), .A(N524), .B(N1025), .CI(N568));
ADDFX1 inst_cellmath__203_0_I689 (.CO(inst_cellmath__203_0_out1[5]), .S(inst_cellmath__203_0_out0[4]), .A(N1380), .B(N596), .CI(N1383));
ADDFX1 inst_cellmath__203_0_I690 (.CO(N1388), .S(N1387), .A(N1027), .B(inst_cellmath__203_0_in0[2]), .CI(N1077));
ADDFX1 inst_cellmath__203_0_I691 (.CO(N1390), .S(N1389), .A(N526), .B(N1387), .CI(N569));
ADDFX1 inst_cellmath__203_0_I692 (.CO(N1392), .S(N1391), .A(N597), .B(N5666), .CI(N625));
ADDFX1 inst_cellmath__203_0_I693 (.CO(inst_cellmath__203_0_out1[6]), .S(inst_cellmath__203_0_out0[5]), .A(N1389), .B(N1384), .CI(N1391));
ADDFX1 inst_cellmath__203_0_I694 (.CO(N1396), .S(N1395), .A(N1078), .B(N1029), .CI(N1388));
ADDFX1 inst_cellmath__203_0_I695 (.CO(N1398), .S(N1397), .A(N528), .B(N1395), .CI(N570));
ADDFX1 inst_cellmath__203_0_I696 (.CO(N1400), .S(N1399), .A(N626), .B(N598), .CI(N1390));
ADDFX1 inst_cellmath__203_0_I697 (.CO(inst_cellmath__203_0_out1[7]), .S(inst_cellmath__203_0_out0[6]), .A(N1392), .B(N1397), .CI(N1399));
ADDFX1 inst_cellmath__203_0_I698 (.CO(N1404), .S(N1403), .A(N1031), .B(N5721), .CI(N1109));
ADDFX1 inst_cellmath__203_0_I699 (.CO(N1406), .S(N1405), .A(N1403), .B(N1079), .CI(N1396));
ADDFX1 inst_cellmath__203_0_I700 (.CO(N1408), .S(N1407), .A(N530), .B(N1405), .CI(N571));
ADDFX1 inst_cellmath__203_0_I701 (.CO(N1410), .S(N1409), .A(N599), .B(N5671), .CI(N627));
ADDFX1 inst_cellmath__203_0_I702 (.CO(N1412), .S(N1411), .A(N1398), .B(N655), .CI(N1407));
ADDFX1 inst_cellmath__203_0_I703 (.CO(inst_cellmath__203_0_out1[8]), .S(inst_cellmath__203_0_out0[7]), .A(N1409), .B(N1400), .CI(N1411));
ADDFX1 inst_cellmath__203_0_I704 (.CO(N1416), .S(N1415), .A(N1110), .B(N1033), .CI(N1080));
ADDFX1 inst_cellmath__203_0_I705 (.CO(N1418), .S(N1417), .A(N1415), .B(N1404), .CI(N1406));
ADDFX1 inst_cellmath__203_0_I706 (.CO(N1420), .S(N1419), .A(N532), .B(N1417), .CI(N572));
ADDFX1 inst_cellmath__203_0_I707 (.CO(N1422), .S(N1421), .A(N628), .B(N600), .CI(N656));
ADDFX1 inst_cellmath__203_0_I708 (.CO(N1424), .S(N1423), .A(N1419), .B(N1408), .CI(N1410));
ADDFX1 inst_cellmath__203_0_I709 (.CO(inst_cellmath__203_0_out1[9]), .S(inst_cellmath__203_0_out0[8]), .A(N1421), .B(N1412), .CI(N1423));
ADDFX1 inst_cellmath__203_0_I710 (.CO(N1428), .S(N1427), .A(N1035), .B(N5726), .CI(N1141));
ADDFX1 inst_cellmath__203_0_I711 (.CO(N1430), .S(N1429), .A(N1081), .B(N1111), .CI(N1416));
ADDFX1 inst_cellmath__203_0_I712 (.CO(N1432), .S(N1431), .A(N1429), .B(N1427), .CI(N1418));
ADDFX1 inst_cellmath__203_0_I713 (.CO(N1434), .S(N1433), .A(N1431), .B(N534), .CI(N5676));
ADDFX1 inst_cellmath__203_0_I714 (.CO(N1436), .S(N1435), .A(N685), .B(N573), .CI(N601));
ADDFX1 inst_cellmath__203_0_I715 (.CO(N1438), .S(N1437), .A(N657), .B(N629), .CI(N1420));
ADDFX1 inst_cellmath__203_0_I716 (.CO(N1440), .S(N1439), .A(N1422), .B(N1433), .CI(N1435));
ADDFX1 inst_cellmath__203_0_I717 (.CO(inst_cellmath__203_0_out1[10]), .S(inst_cellmath__203_0_out0[9]), .A(N1424), .B(N1437), .CI(N1439));
ADDFX1 inst_cellmath__203_0_I718 (.CO(N1444), .S(N1443), .A(N1142), .B(N1037), .CI(N1112));
ADDFX1 inst_cellmath__203_0_I719 (.CO(N1446), .S(N1445), .A(N1428), .B(N1082), .CI(N1443));
ADDFX1 inst_cellmath__203_0_I720 (.CO(N1448), .S(N1447), .A(N1445), .B(N1430), .CI(N1432));
ADDFX1 inst_cellmath__203_0_I721 (.CO(N1450), .S(N1449), .A(N1447), .B(N536), .CI(N574));
ADDFX1 inst_cellmath__203_0_I722 (.CO(N1452), .S(N1451), .A(N602), .B(N686), .CI(N630));
ADDFX1 inst_cellmath__203_0_I723 (.CO(N1454), .S(N1453), .A(N1434), .B(N658), .CI(N1449));
ADDFX1 inst_cellmath__203_0_I724 (.CO(N1456), .S(N1455), .A(N1438), .B(N1436), .CI(N1451));
ADDFX1 inst_cellmath__203_0_I725 (.CO(inst_cellmath__203_0_out1[11]), .S(inst_cellmath__203_0_out0[10]), .A(N1440), .B(N1453), .CI(N1455));
ADDFX1 inst_cellmath__203_0_I726 (.CO(N1460), .S(N1459), .A(N1039), .B(N5731), .CI(N1173));
ADDFX1 inst_cellmath__203_0_I727 (.CO(N1462), .S(N1461), .A(N1113), .B(N1143), .CI(N1083));
ADDFX1 inst_cellmath__203_0_I728 (.CO(N1464), .S(N1463), .A(N1459), .B(N1444), .CI(N1461));
ADDFX1 inst_cellmath__203_0_I729 (.CO(N1466), .S(N1465), .A(N1463), .B(N1446), .CI(N538));
ADDFX1 inst_cellmath__203_0_I730 (.CO(N1468), .S(N1467), .A(N1465), .B(N1448), .CI(N575));
ADDFX1 inst_cellmath__203_0_I731 (.CO(N1470), .S(N1469), .A(N687), .B(N5681), .CI(N603));
ADDFX1 inst_cellmath__203_0_I732 (.CO(N1472), .S(N1471), .A(N715), .B(N631), .CI(N659));
ADDFX1 inst_cellmath__203_0_I733 (.CO(N1474), .S(N1473), .A(N1467), .B(N1450), .CI(N1452));
ADDFX1 inst_cellmath__203_0_I734 (.CO(N1476), .S(N1475), .A(N1454), .B(N1469), .CI(N1471));
ADDFX1 inst_cellmath__203_0_I735 (.CO(inst_cellmath__203_0_out1[12]), .S(inst_cellmath__203_0_out0[11]), .A(N1456), .B(N1473), .CI(N1475));
ADDFX1 inst_cellmath__203_0_I736 (.CO(N1480), .S(N1479), .A(N1174), .B(N1041), .CI(N1144));
ADDFX1 inst_cellmath__203_0_I737 (.CO(N1482), .S(N1481), .A(N1084), .B(N1114), .CI(N1460));
ADDFX1 inst_cellmath__203_0_I738 (.CO(N1484), .S(N1483), .A(N1479), .B(N1462), .CI(N1481));
ADDFX1 inst_cellmath__203_0_I739 (.CO(N1486), .S(N1485), .A(N1483), .B(N1464), .CI(N540));
ADDFX1 inst_cellmath__203_0_I740 (.CO(N1488), .S(N1487), .A(N1485), .B(N1466), .CI(N576));
ADDFX1 inst_cellmath__203_0_I741 (.CO(N1490), .S(N1489), .A(N604), .B(N688), .CI(N632));
ADDFX1 inst_cellmath__203_0_I742 (.CO(N1492), .S(N1491), .A(N716), .B(N660), .CI(N1468));
ADDFX1 inst_cellmath__203_0_I743 (.CO(N1494), .S(N1493), .A(N1470), .B(N1487), .CI(N1472));
ADDFX1 inst_cellmath__203_0_I744 (.CO(N1496), .S(N1495), .A(N1491), .B(N1489), .CI(N1474));
ADDFX1 inst_cellmath__203_0_I745 (.CO(inst_cellmath__203_0_out1[13]), .S(inst_cellmath__203_0_out0[12]), .A(N1476), .B(N1493), .CI(N1495));
ADDFX1 inst_cellmath__203_0_I746 (.CO(N1500), .S(N1499), .A(N1043), .B(N5736), .CI(N1205));
ADDFX1 inst_cellmath__203_0_I747 (.CO(N1502), .S(N1501), .A(N1085), .B(N1175), .CI(N1145));
ADDFX1 inst_cellmath__203_0_I748 (.CO(N1504), .S(N1503), .A(N1480), .B(N1115), .CI(N1499));
ADDFX1 inst_cellmath__203_0_I749 (.CO(N1506), .S(N1505), .A(N1501), .B(N1482), .CI(N1503));
ADDFX1 inst_cellmath__203_0_I750 (.CO(N1508), .S(N1507), .A(N1505), .B(N1484), .CI(N542));
ADDFX1 inst_cellmath__203_0_I751 (.CO(N1510), .S(N1509), .A(N1507), .B(N1486), .CI(N577));
ADDFX1 inst_cellmath__203_0_I752 (.CO(N1512), .S(N1511), .A(N5686), .B(N689), .CI(N717));
ADDFX1 inst_cellmath__203_0_I753 (.CO(N1514), .S(N1513), .A(N633), .B(N605), .CI(N661));
ADDFX1 inst_cellmath__203_0_I754 (.CO(N1516), .S(N1515), .A(N1488), .B(N745), .CI(N1509));
ADDFX1 inst_cellmath__203_0_I755 (.CO(N1518), .S(N1517), .A(N1492), .B(N1490), .CI(N1511));
ADDFX1 inst_cellmath__203_0_I756 (.CO(N1520), .S(N1519), .A(N1494), .B(N1513), .CI(N1515));
ADDFX1 inst_cellmath__203_0_I757 (.CO(inst_cellmath__203_0_out1[14]), .S(inst_cellmath__203_0_out0[13]), .A(N1517), .B(N1496), .CI(N1519));
ADDFX1 inst_cellmath__203_0_I758 (.CO(N1524), .S(N1523), .A(N1206), .B(N1045), .CI(N1176));
ADDFX1 inst_cellmath__203_0_I759 (.CO(N1526), .S(N1525), .A(N1086), .B(N1146), .CI(N1116));
ADDFX1 inst_cellmath__203_0_I760 (.CO(N1528), .S(N1527), .A(N1502), .B(N1500), .CI(N1523));
ADDFX1 inst_cellmath__203_0_I761 (.CO(N1530), .S(N1529), .A(N1504), .B(N1525), .CI(N1527));
ADDFX1 inst_cellmath__203_0_I762 (.CO(N1532), .S(N1531), .A(N1529), .B(N1506), .CI(N544));
ADDFX1 inst_cellmath__203_0_I763 (.CO(N1534), .S(N1533), .A(N1531), .B(N1508), .CI(N578));
ADDFX1 inst_cellmath__203_0_I764 (.CO(N1536), .S(N1535), .A(N606), .B(N690), .CI(N634));
ADDFX1 inst_cellmath__203_0_I765 (.CO(N1538), .S(N1537), .A(N718), .B(N662), .CI(N746));
ADDFX1 inst_cellmath__203_0_I766 (.CO(N1540), .S(N1539), .A(N1533), .B(N1510), .CI(N1512));
ADDFX1 inst_cellmath__203_0_I767 (.CO(N1542), .S(N1541), .A(N1535), .B(N1514), .CI(N1516));
ADDFX1 inst_cellmath__203_0_I768 (.CO(N1544), .S(N1543), .A(N1539), .B(N1537), .CI(N1518));
ADDFX1 inst_cellmath__203_0_I769 (.CO(inst_cellmath__203_0_out1[15]), .S(inst_cellmath__203_0_out0[14]), .A(N1520), .B(N1541), .CI(N1543));
ADDHX1 inst_cellmath__203_0_I770 (.CO(N1548), .S(N1547), .A(N5741), .B(N1047));
ADDFX1 inst_cellmath__203_0_I771 (.CO(N1550), .S(N1549), .A(N1547), .B(N1237), .CI(N1207));
ADDFX1 inst_cellmath__203_0_I772 (.CO(N1552), .S(N1551), .A(N1177), .B(N1117), .CI(N1147));
ADDFX1 inst_cellmath__203_0_I773 (.CO(N1554), .S(N1553), .A(N1524), .B(N1087), .CI(N1526));
ADDFX1 inst_cellmath__203_0_I774 (.CO(N1556), .S(N1555), .A(N1551), .B(N1549), .CI(N1528));
ADDFX1 inst_cellmath__203_0_I775 (.CO(N1558), .S(N1557), .A(N1555), .B(N1553), .CI(N1530));
ADDFX1 inst_cellmath__203_0_I776 (.CO(N1560), .S(N1559), .A(N1557), .B(N546), .CI(N1532));
ADDFX1 inst_cellmath__203_0_I777 (.CO(N1562), .S(N1561), .A(N779), .B(N1559), .CI(N579));
ADDFX1 inst_cellmath__203_0_I778 (.CO(N1564), .S(N1563), .A(N607), .B(N691), .CI(N635));
ADDFX1 inst_cellmath__203_0_I779 (.CO(N1566), .S(N1565), .A(N719), .B(N663), .CI(N747));
ADDFX1 inst_cellmath__203_0_I780 (.CO(N1568), .S(N1567), .A(N1561), .B(N1534), .CI(N1536));
ADDFX1 inst_cellmath__203_0_I781 (.CO(N1570), .S(N1569), .A(N1563), .B(N1538), .CI(N1565));
ADDFX1 inst_cellmath__203_0_I782 (.CO(N1572), .S(N1571), .A(N1567), .B(N1540), .CI(N1542));
ADDFX1 inst_cellmath__203_0_I783 (.CO(inst_cellmath__203_0_out1[16]), .S(inst_cellmath__203_0_out0[15]), .A(N1569), .B(N1544), .CI(N1571));
ADDFX1 inst_cellmath__203_0_I784 (.CO(N1576), .S(N1575), .A(N1548), .B(N1049), .CI(N1238));
ADDFX1 inst_cellmath__203_0_I785 (.CO(N1578), .S(N1577), .A(N1178), .B(N1208), .CI(N1148));
ADDFX1 inst_cellmath__203_0_I786 (.CO(N1580), .S(N1579), .A(N1088), .B(N1118), .CI(N1550));
ADDFX1 inst_cellmath__203_0_I787 (.CO(N1582), .S(N1581), .A(N1575), .B(N1552), .CI(N1577));
ADDFX1 inst_cellmath__203_0_I788 (.CO(N1584), .S(N1583), .A(N1579), .B(N1554), .CI(N1581));
ADDFX1 inst_cellmath__203_0_I789 (.CO(N1586), .S(N1585), .A(N548), .B(N1556), .CI(N1583));
ADDFX1 inst_cellmath__203_0_I790 (.CO(N1588), .S(N1587), .A(N1585), .B(N1558), .CI(N1560));
ADDFX1 inst_cellmath__203_0_I791 (.CO(N1590), .S(N1589), .A(N1587), .B(N781), .CI(N580));
ADDFX1 inst_cellmath__203_0_I792 (.CO(N1592), .S(N1591), .A(N608), .B(N692), .CI(N636));
ADDFX1 inst_cellmath__203_0_I793 (.CO(N1594), .S(N1593), .A(N720), .B(N664), .CI(N748));
ADDFX1 inst_cellmath__203_0_I794 (.CO(N1596), .S(N1595), .A(N1589), .B(N1562), .CI(N1564));
ADDFX1 inst_cellmath__203_0_I795 (.CO(N1598), .S(N1597), .A(N1591), .B(N1566), .CI(N1593));
ADDFX1 inst_cellmath__203_0_I796 (.CO(N1600), .S(N1599), .A(N1595), .B(N1568), .CI(N1570));
ADDFX1 inst_cellmath__203_0_I797 (.CO(inst_cellmath__203_0_out1[17]), .S(inst_cellmath__203_0_out0[16]), .A(N1572), .B(N1597), .CI(N1599));
ADDFX1 inst_cellmath__203_0_I798 (.CO(N1604), .S(N1603), .A(N1051), .B(N5746), .CI(N1269));
ADDFX1 inst_cellmath__203_0_I799 (.CO(N1606), .S(N1605), .A(N1149), .B(N1089), .CI(N1239));
ADDFX1 inst_cellmath__203_0_I800 (.CO(N1608), .S(N1607), .A(N1179), .B(N1209), .CI(N1119));
ADDFX1 inst_cellmath__203_0_I801 (.CO(N1610), .S(N1609), .A(N1578), .B(N1576), .CI(N1603));
ADDFX1 inst_cellmath__203_0_I802 (.CO(N1612), .S(N1611), .A(N1580), .B(N1605), .CI(N1607));
ADDFX1 inst_cellmath__203_0_I803 (.CO(N1614), .S(N1613), .A(N1609), .B(N1582), .CI(N1611));
ADDFX1 inst_cellmath__203_0_I804 (.CO(N1616), .S(N1615), .A(N550), .B(N1584), .CI(N1613));
ADDFX1 inst_cellmath__203_0_I805 (.CO(N1618), .S(N1617), .A(N1615), .B(N1586), .CI(N1588));
ADDFX1 inst_cellmath__203_0_I806 (.CO(N1620), .S(N1619), .A(N581), .B(N783), .CI(N693));
ADDFX1 inst_cellmath__203_0_I807 (.CO(N1622), .S(N1621), .A(N1617), .B(N609), .CI(N721));
ADDFX1 inst_cellmath__203_0_I808 (.CO(N1624), .S(N1623), .A(N665), .B(N637), .CI(N749));
ADDFX1 inst_cellmath__203_0_I809 (.CO(N1626), .S(N1625), .A(N1592), .B(N1590), .CI(N1619));
ADDFX1 inst_cellmath__203_0_I810 (.CO(N1628), .S(N1627), .A(N1621), .B(N1594), .CI(N1623));
ADDFX1 inst_cellmath__203_0_I811 (.CO(N1630), .S(N1629), .A(N1625), .B(N1596), .CI(N1598));
ADDFX1 inst_cellmath__203_0_I812 (.CO(inst_cellmath__203_0_out1[18]), .S(inst_cellmath__203_0_out0[17]), .A(N1600), .B(N1627), .CI(N1629));
ADDFX1 inst_cellmath__203_0_I813 (.CO(N1634), .S(N1633), .A(N1270), .B(N1053), .CI(N1240));
ADDFX1 inst_cellmath__203_0_I814 (.CO(N1636), .S(N1635), .A(N1210), .B(N1090), .CI(N1180));
ADDFX1 inst_cellmath__203_0_I815 (.CO(N1638), .S(N1637), .A(N1120), .B(N1150), .CI(N1604));
ADDFX1 inst_cellmath__203_0_I816 (.CO(N1640), .S(N1639), .A(N1608), .B(N1606), .CI(N1633));
ADDFX1 inst_cellmath__203_0_I817 (.CO(N1642), .S(N1641), .A(N1637), .B(N1635), .CI(N1610));
ADDFX1 inst_cellmath__203_0_I818 (.CO(N1644), .S(N1643), .A(N1639), .B(N1612), .CI(N1641));
ADDFX1 inst_cellmath__203_0_I819 (.CO(N1646), .S(N1645), .A(N552), .B(N1614), .CI(N1643));
ADDFX1 inst_cellmath__203_0_I820 (.CO(N1648), .S(N1647), .A(N1645), .B(N1616), .CI(N785));
ADDFX1 inst_cellmath__203_0_I821 (.CO(N1650), .S(N1649), .A(N582), .B(N1618), .CI(N694));
ADDFX1 inst_cellmath__203_0_I822 (.CO(N1652), .S(N1651), .A(N638), .B(N610), .CI(N722));
ADDFX1 inst_cellmath__203_0_I823 (.CO(N1654), .S(N1653), .A(N1647), .B(N666), .CI(N750));
ADDFX1 inst_cellmath__203_0_I824 (.CO(N1656), .S(N1655), .A(N1622), .B(N1620), .CI(N1649));
ADDFX1 inst_cellmath__203_0_I825 (.CO(N1658), .S(N1657), .A(N1651), .B(N1624), .CI(N1653));
ADDFX1 inst_cellmath__203_0_I826 (.CO(N1660), .S(N1659), .A(N1655), .B(N1626), .CI(N1628));
ADDFX1 inst_cellmath__203_0_I827 (.CO(inst_cellmath__203_0_out1[19]), .S(inst_cellmath__203_0_out0[18]), .A(N1630), .B(N1657), .CI(N1659));
ADDFX1 inst_cellmath__203_0_I828 (.CO(N1664), .S(N1663), .A(N1055), .B(N5751), .CI(N1301));
ADDFX1 inst_cellmath__203_0_I829 (.CO(N1666), .S(N1665), .A(N1181), .B(N1121), .CI(N1271));
ADDFX1 inst_cellmath__203_0_I830 (.CO(N1668), .S(N1667), .A(N1241), .B(N1091), .CI(N1211));
ADDFX1 inst_cellmath__203_0_I831 (.CO(N1670), .S(N1669), .A(N1634), .B(N1151), .CI(N1636));
ADDFX1 inst_cellmath__203_0_I832 (.CO(N1672), .S(N1671), .A(N1638), .B(N1663), .CI(N1665));
ADDFX1 inst_cellmath__203_0_I833 (.CO(N1674), .S(N1673), .A(N1640), .B(N1667), .CI(N1669));
ADDFX1 inst_cellmath__203_0_I834 (.CO(N1676), .S(N1675), .A(N1642), .B(N1671), .CI(N1673));
ADDFX1 inst_cellmath__203_0_I835 (.CO(N1678), .S(N1677), .A(N1644), .B(N554), .CI(N1675));
ADDFX1 inst_cellmath__203_0_I836 (.CO(N1680), .S(N1679), .A(N1677), .B(N1646), .CI(N787));
ADDFX1 inst_cellmath__203_0_I837 (.CO(N1682), .S(N1681), .A(N1648), .B(N583), .CI(N695));
ADDFX1 inst_cellmath__203_0_I838 (.CO(N1684), .S(N1683), .A(N639), .B(N611), .CI(N723));
ADDFX1 inst_cellmath__203_0_I839 (.CO(N1686), .S(N1685), .A(N1679), .B(N667), .CI(N751));
ADDFX1 inst_cellmath__203_0_I840 (.CO(N1688), .S(N1687), .A(N1652), .B(N1650), .CI(N1681));
ADDFX1 inst_cellmath__203_0_I841 (.CO(N1690), .S(N1689), .A(N1683), .B(N1654), .CI(N1685));
ADDFX1 inst_cellmath__203_0_I842 (.CO(N1692), .S(N1691), .A(N1687), .B(N1656), .CI(N1658));
ADDFX1 inst_cellmath__203_0_I843 (.CO(inst_cellmath__203_0_out1[20]), .S(inst_cellmath__203_0_out0[19]), .A(N1660), .B(N1689), .CI(N1691));
INVXL fap1_A_I1798 (.Y(N5461), .A(N1732));
ADDFX1 fap1_A_I1799 (.CO(N1696), .S(N1695), .A(N1272), .B(N1302), .CI(N5461));
ADDFX1 inst_cellmath__203_0_I845 (.CO(N1700), .S(N1699), .A(N1092), .B(N1122), .CI(N1242));
ADDFX1 inst_cellmath__203_0_I846 (.CO(N1702), .S(N1701), .A(N1212), .B(N1182), .CI(N1152));
ADDFX1 inst_cellmath__203_0_I847 (.CO(N1704), .S(N1703), .A(N1666), .B(N1664), .CI(N1668));
ADDFX1 inst_cellmath__203_0_I848 (.CO(N1706), .S(N1705), .A(N1699), .B(N1695), .CI(N1701));
ADDFX1 inst_cellmath__203_0_I849 (.CO(N1708), .S(N1707), .A(N1672), .B(N1670), .CI(N1703));
ADDFX1 inst_cellmath__203_0_I850 (.CO(N1710), .S(N1709), .A(N1674), .B(N1705), .CI(N1707));
ADDFX1 inst_cellmath__203_0_I851 (.CO(N1712), .S(N1711), .A(N1676), .B(N5655), .CI(N1709));
ADDFX1 inst_cellmath__203_0_I852 (.CO(N1714), .S(N1713), .A(N1711), .B(N1678), .CI(N789));
ADDFX1 inst_cellmath__203_0_I853 (.CO(N1716), .S(N1715), .A(N1680), .B(N584), .CI(N696));
ADDFX1 inst_cellmath__203_0_I854 (.CO(N1718), .S(N1717), .A(N640), .B(N612), .CI(N724));
ADDFX1 inst_cellmath__203_0_I855 (.CO(N1720), .S(N1719), .A(N1713), .B(N668), .CI(N752));
ADDFX1 inst_cellmath__203_0_I856 (.CO(N1722), .S(N1721), .A(N1684), .B(N1682), .CI(N1715));
ADDFX1 inst_cellmath__203_0_I857 (.CO(N1724), .S(N1723), .A(N1717), .B(N1686), .CI(N1719));
ADDFX1 inst_cellmath__203_0_I858 (.CO(N1726), .S(N1725), .A(N1721), .B(N1688), .CI(N1690));
ADDFX1 inst_cellmath__203_0_I859 (.CO(inst_cellmath__203_0_out1[21]), .S(inst_cellmath__203_0_out0[20]), .A(N1692), .B(N1723), .CI(N1725));
ADDFX1 inst_cellmath__203_0_I1801 (.CO(N1730), .S(N1729), .A(N1093), .B(N1059), .CI(N5461));
ADDFX1 inst_cellmath__203_0_I861 (.CO(N1734), .S(N1733), .A(N1213), .B(N1153), .CI(N1303));
ADDFX1 inst_cellmath__203_0_I862 (.CO(N1736), .S(N1735), .A(N1273), .B(N1123), .CI(N1243));
ADDFX1 inst_cellmath__203_0_I863 (.CO(N1738), .S(N1737), .A(N1696), .B(N1183), .CI(N1700));
ADDFX1 inst_cellmath__203_0_I864 (.CO(N1740), .S(N1739), .A(N1729), .B(N1702), .CI(N1733));
ADDFX1 inst_cellmath__203_0_I865 (.CO(N1742), .S(N1741), .A(N1704), .B(N1735), .CI(N1737));
ADDFX1 inst_cellmath__203_0_I866 (.CO(N1744), .S(N1743), .A(N1739), .B(N1706), .CI(N1708));
ADDFX1 inst_cellmath__203_0_I867 (.CO(N1746), .S(N1745), .A(N1710), .B(N1741), .CI(N1743));
ADDFX1 inst_cellmath__203_0_I868 (.CO(N1748), .S(N1747), .A(N1745), .B(N1712), .CI(N791));
ADDFX1 inst_cellmath__203_0_I869 (.CO(N1750), .S(N1749), .A(N1714), .B(N585), .CI(N697));
ADDFX1 inst_cellmath__203_0_I870 (.CO(N1752), .S(N1751), .A(N641), .B(N613), .CI(N725));
ADDFX1 inst_cellmath__203_0_I871 (.CO(N1754), .S(N1753), .A(N1747), .B(N669), .CI(N753));
ADDFX1 inst_cellmath__203_0_I872 (.CO(N1756), .S(N1755), .A(N1718), .B(N1716), .CI(N1749));
ADDFX1 inst_cellmath__203_0_I873 (.CO(N1758), .S(N1757), .A(N1751), .B(N1720), .CI(N1753));
ADDFX1 inst_cellmath__203_0_I874 (.CO(N1760), .S(N1759), .A(N1755), .B(N1722), .CI(N1724));
ADDFX1 inst_cellmath__203_0_I875 (.CO(inst_cellmath__203_0_out1[22]), .S(inst_cellmath__203_0_out0[21]), .A(N1726), .B(N1757), .CI(N1759));
ADDFX1 inst_cellmath__203_0_I876 (.CO(N1764), .S(N1763), .A(N1061), .B(N1732), .CI(N1154));
ADDFX1 inst_cellmath__203_0_I877 (.CO(N1766), .S(N1765), .A(N1304), .B(N1124), .CI(N1274));
ADDFX1 inst_cellmath__203_0_I878 (.CO(N1768), .S(N1767), .A(N1244), .B(N1214), .CI(N1184));
ADDFX1 inst_cellmath__203_0_I879 (.CO(N1770), .S(N1769), .A(N1730), .B(N1094), .CI(N1734));
ADDFX1 inst_cellmath__203_0_I880 (.CO(N1772), .S(N1771), .A(N1763), .B(N1736), .CI(N1765));
ADDFX1 inst_cellmath__203_0_I881 (.CO(N1774), .S(N1773), .A(N1738), .B(N1767), .CI(N1769));
ADDFX1 inst_cellmath__203_0_I882 (.CO(N1776), .S(N1775), .A(N1771), .B(N1740), .CI(N1742));
ADDFX1 inst_cellmath__203_0_I883 (.CO(N1778), .S(N1777), .A(N1744), .B(N1773), .CI(N1775));
ADDFX1 inst_cellmath__203_0_I884 (.CO(N1780), .S(N1779), .A(N1777), .B(N1746), .CI(N5659));
ADDFX1 inst_cellmath__203_0_I885 (.CO(N1782), .S(N1781), .A(N1748), .B(N793), .CI(N1779));
ADDFX1 inst_cellmath__203_0_I886 (.CO(N1784), .S(N1783), .A(N614), .B(N698), .CI(N642));
ADDFX1 inst_cellmath__203_0_I887 (.CO(N1786), .S(N1785), .A(N726), .B(N670), .CI(N754));
ADDFX1 inst_cellmath__203_0_I888 (.CO(N1788), .S(N1787), .A(N1781), .B(N1750), .CI(N1752));
ADDFX1 inst_cellmath__203_0_I889 (.CO(N1790), .S(N1789), .A(N1783), .B(N1754), .CI(N1785));
ADDFX1 inst_cellmath__203_0_I890 (.CO(N1792), .S(N1791), .A(N1787), .B(N1756), .CI(N1758));
ADDFX1 inst_cellmath__203_0_I891 (.CO(inst_cellmath__203_0_out1[23]), .S(inst_cellmath__203_0_out0[22]), .A(N1760), .B(N1789), .CI(N1791));
INVXL fap1_A_I1802 (.Y(N5479), .A(N1798));
ADDFX1 fap1_A_I1803 (.CO(N1796), .S(N1795), .A(N1185), .B(N1125), .CI(N5479));
ADDFX1 inst_cellmath__203_0_I893 (.CO(N1800), .S(N1799), .A(N1245), .B(N1155), .CI(N1305));
ADDFX1 inst_cellmath__203_0_I894 (.CO(N1802), .S(N1801), .A(N1275), .B(N1095), .CI(N1215));
ADDFX1 inst_cellmath__203_0_I895 (.CO(N1804), .S(N1803), .A(N1766), .B(N1764), .CI(N1768));
ADDFX1 inst_cellmath__203_0_I896 (.CO(N1806), .S(N1805), .A(N1799), .B(N1795), .CI(N1801));
ADDFX1 inst_cellmath__203_0_I897 (.CO(N1808), .S(N1807), .A(N1772), .B(N1770), .CI(N1803));
ADDFX1 inst_cellmath__203_0_I898 (.CO(N1810), .S(N1809), .A(N1774), .B(N1805), .CI(N1807));
ADDFX1 inst_cellmath__203_0_I899 (.CO(N1812), .S(N1811), .A(N1809), .B(N1776), .CI(N1778));
ADDFX1 inst_cellmath__203_0_I900 (.CO(N1814), .S(N1813), .A(N795), .B(N1811), .CI(N1780));
ADDFX1 inst_cellmath__203_0_I901 (.CO(N1816), .S(N1815), .A(N615), .B(N699), .CI(N643));
ADDFX1 inst_cellmath__203_0_I902 (.CO(N1818), .S(N1817), .A(N727), .B(N671), .CI(N755));
ADDFX1 inst_cellmath__203_0_I903 (.CO(N1820), .S(N1819), .A(N1782), .B(N1813), .CI(N1784));
ADDFX1 inst_cellmath__203_0_I904 (.CO(N1822), .S(N1821), .A(N1815), .B(N1786), .CI(N1817));
ADDFX1 inst_cellmath__203_0_I905 (.CO(N1824), .S(N1823), .A(N1819), .B(N1788), .CI(N1790));
ADDFX1 inst_cellmath__203_0_I906 (.CO(inst_cellmath__203_0_out1[24]), .S(inst_cellmath__203_0_out0[23]), .A(N1792), .B(N1821), .CI(N1823));
INVXL fap1_A_I1804 (.Y(N5488), .A(N1830));
ADDFX1 fap1_A_I1805 (.CO(N1828), .S(N1827), .A(N1186), .B(N1798), .CI(N5488));
ADDFX1 inst_cellmath__203_0_I908 (.CO(N1832), .S(N1831), .A(N1306), .B(N1156), .CI(N1126));
ADDFX1 inst_cellmath__203_0_I909 (.CO(N1834), .S(N1833), .A(N1246), .B(N1096), .CI(N1276));
ADDFX1 inst_cellmath__203_0_I910 (.CO(N1836), .S(N1835), .A(N1796), .B(N1216), .CI(N1800));
ADDFX1 inst_cellmath__203_0_I911 (.CO(N1838), .S(N1837), .A(N1827), .B(N1802), .CI(N1831));
ADDFX1 inst_cellmath__203_0_I912 (.CO(N1840), .S(N1839), .A(N1804), .B(N1833), .CI(N1835));
ADDFX1 inst_cellmath__203_0_I913 (.CO(N1842), .S(N1841), .A(N1837), .B(N1806), .CI(N1808));
ADDFX1 inst_cellmath__203_0_I914 (.CO(N1844), .S(N1843), .A(N1810), .B(N1839), .CI(N1841));
ADDFX1 inst_cellmath__203_0_I915 (.CO(N1846), .S(N1845), .A(N1812), .B(N1843), .CI(N5664));
ADDFX1 inst_cellmath__203_0_I916 (.CO(N1848), .S(N1847), .A(N1845), .B(N797), .CI(N700));
ADDFX1 inst_cellmath__203_0_I917 (.CO(N1850), .S(N1849), .A(N728), .B(N1814), .CI(N672));
ADDFX1 inst_cellmath__203_0_I918 (.CO(N1852), .S(N1851), .A(N756), .B(N644), .CI(N1816));
ADDFX1 inst_cellmath__203_0_I919 (.CO(N1854), .S(N1853), .A(N1818), .B(N1847), .CI(N1849));
ADDFX1 inst_cellmath__203_0_I920 (.CO(N1856), .S(N1855), .A(N1851), .B(N1820), .CI(N1822));
ADDFX1 inst_cellmath__203_0_I921 (.CO(inst_cellmath__203_0_out1[25]), .S(inst_cellmath__203_0_out0[24]), .A(N1824), .B(N1853), .CI(N1855));
XNOR2X1 hap1_A_I1806 (.Y(N1859), .A(N1067), .B(N1830));
OR2XL hap1_A_I1807 (.Y(N1860), .A(N1067), .B(N1830));
ADDFX1 inst_cellmath__203_0_I923 (.CO(N1864), .S(N1863), .A(N1157), .B(N1859), .CI(N1277));
ADDFX1 inst_cellmath__203_0_I924 (.CO(N1866), .S(N1865), .A(N1187), .B(N1217), .CI(N1097));
ADDFX1 inst_cellmath__203_0_I925 (.CO(N1868), .S(N1867), .A(N1307), .B(N1127), .CI(N1247));
ADDFX1 inst_cellmath__203_0_I926 (.CO(N1870), .S(N1869), .A(N1832), .B(N1828), .CI(N1834));
ADDFX1 inst_cellmath__203_0_I927 (.CO(N1872), .S(N1871), .A(N1865), .B(N1863), .CI(N1867));
ADDFX1 inst_cellmath__203_0_I928 (.CO(N1874), .S(N1873), .A(N1838), .B(N1836), .CI(N1869));
ADDFX1 inst_cellmath__203_0_I929 (.CO(N1876), .S(N1875), .A(N1840), .B(N1871), .CI(N1873));
ADDFX1 inst_cellmath__203_0_I930 (.CO(N1878), .S(N1877), .A(N1875), .B(N1842), .CI(N1844));
ADDFX1 inst_cellmath__203_0_I931 (.CO(N1880), .S(N1879), .A(N1877), .B(N799), .CI(N1846));
ADDFX1 inst_cellmath__203_0_I932 (.CO(N1882), .S(N1881), .A(N645), .B(N701), .CI(N729));
ADDFX1 inst_cellmath__203_0_I933 (.CO(N1884), .S(N1883), .A(N757), .B(N673), .CI(N1879));
ADDFX1 inst_cellmath__203_0_I934 (.CO(N1886), .S(N1885), .A(N1850), .B(N1848), .CI(N1881));
ADDFX1 inst_cellmath__203_0_I935 (.CO(N1888), .S(N1887), .A(N1883), .B(N1852), .CI(N1854));
ADDFX1 inst_cellmath__203_0_I936 (.CO(inst_cellmath__203_0_out1[26]), .S(inst_cellmath__203_0_out0[25]), .A(N1856), .B(N1885), .CI(N1887));
ADDHX1 inst_cellmath__203_0_I937 (.CO(N1892), .S(N1891), .A(N1860), .B(N1098));
ADDFX1 inst_cellmath__203_0_I938 (.CO(N1894), .S(N1893), .A(N1218), .B(N1891), .CI(N1188));
ADDFX1 inst_cellmath__203_0_I939 (.CO(N1896), .S(N1895), .A(N1278), .B(N1128), .CI(N1308));
ADDFX1 inst_cellmath__203_0_I940 (.CO(N1898), .S(N1897), .A(N1248), .B(N1158), .CI(N1864));
ADDFX1 inst_cellmath__203_0_I941 (.CO(N1900), .S(N1899), .A(N1868), .B(N1866), .CI(N1893));
ADDFX1 inst_cellmath__203_0_I942 (.CO(N1902), .S(N1901), .A(N1870), .B(N1895), .CI(N1897));
ADDFX1 inst_cellmath__203_0_I943 (.CO(N1904), .S(N1903), .A(N1899), .B(N1872), .CI(N1874));
ADDFX1 inst_cellmath__203_0_I944 (.CO(N1906), .S(N1905), .A(N1903), .B(N1901), .CI(N1876));
ADDFX1 inst_cellmath__203_0_I945 (.CO(N1908), .S(N1907), .A(N1878), .B(N1905), .CI(N5669));
ADDFX1 inst_cellmath__203_0_I946 (.CO(N1910), .S(N1909), .A(N1907), .B(N801), .CI(N702));
ADDFX1 inst_cellmath__203_0_I947 (.CO(N1912), .S(N1911), .A(N730), .B(N674), .CI(N1880));
ADDFX1 inst_cellmath__203_0_I948 (.CO(N1914), .S(N1913), .A(N1882), .B(N758), .CI(N1909));
ADDFX1 inst_cellmath__203_0_I949 (.CO(N1916), .S(N1915), .A(N1911), .B(N1884), .CI(N1886));
ADDFX1 inst_cellmath__203_0_I950 (.CO(inst_cellmath__203_0_out1[27]), .S(inst_cellmath__203_0_out0[26]), .A(N1888), .B(N1913), .CI(N1915));
XNOR2X1 hap1_A_I1808 (.Y(N1919), .A(N1099), .B(N1892));
OR2XL hap1_A_I1809 (.Y(N1920), .A(N1099), .B(N1892));
ADDFX1 inst_cellmath__203_0_I952 (.CO(N1924), .S(N1923), .A(N1189), .B(N1919), .CI(N1309));
ADDFX1 inst_cellmath__203_0_I953 (.CO(N1926), .S(N1925), .A(N1219), .B(N1249), .CI(N1129));
ADDFX1 inst_cellmath__203_0_I954 (.CO(N1928), .S(N1927), .A(N1279), .B(N1159), .CI(N1894));
ADDFX1 inst_cellmath__203_0_I955 (.CO(N1930), .S(N1929), .A(N1923), .B(N1896), .CI(N1925));
ADDFX1 inst_cellmath__203_0_I956 (.CO(N1932), .S(N1931), .A(N1900), .B(N1898), .CI(N1927));
ADDFX1 inst_cellmath__203_0_I957 (.CO(N1934), .S(N1933), .A(N1902), .B(N1929), .CI(N1931));
ADDFX1 inst_cellmath__203_0_I958 (.CO(N1936), .S(N1935), .A(N1933), .B(N1904), .CI(N1906));
ADDFX1 inst_cellmath__203_0_I959 (.CO(N1938), .S(N1937), .A(N1935), .B(N803), .CI(N1908));
ADDFX1 inst_cellmath__203_0_I960 (.CO(N1940), .S(N1939), .A(N675), .B(N703), .CI(N731));
ADDFX1 inst_cellmath__203_0_I961 (.CO(N1942), .S(N1941), .A(N1937), .B(N759), .CI(N1910));
ADDFX1 inst_cellmath__203_0_I962 (.CO(N1944), .S(N1943), .A(N1939), .B(N1912), .CI(N1941));
ADDFX1 inst_cellmath__203_0_I963 (.CO(inst_cellmath__203_0_out1[28]), .S(inst_cellmath__203_0_out0[27]), .A(N1916), .B(N1914), .CI(N1943));
INVXL fap1_A_I1810 (.Y(N5509), .A(N5720));
ADDFX1 fap1_A_I1811 (.CO(N1948), .S(N1947), .A(N1920), .B(N1130), .CI(N5509));
ADDFX1 inst_cellmath__203_0_I965 (.CO(N1952), .S(N1951), .A(N1220), .B(N1250), .CI(N1160));
ADDFX1 inst_cellmath__203_0_I966 (.CO(N1954), .S(N1953), .A(N1190), .B(N1310), .CI(N1280));
ADDFX1 inst_cellmath__203_0_I967 (.CO(N1956), .S(N1955), .A(N1924), .B(N1947), .CI(N1926));
ADDFX1 inst_cellmath__203_0_I968 (.CO(N1958), .S(N1957), .A(N1928), .B(N1951), .CI(N1953));
ADDFX1 inst_cellmath__203_0_I969 (.CO(N1960), .S(N1959), .A(N1930), .B(N1955), .CI(N1957));
ADDFX1 inst_cellmath__203_0_I970 (.CO(N1962), .S(N1961), .A(N1959), .B(N1932), .CI(N1934));
ADDFX1 inst_cellmath__203_0_I971 (.CO(N1964), .S(N1963), .A(N1936), .B(N1961), .CI(N5674));
ADDFX1 inst_cellmath__203_0_I972 (.CO(N1966), .S(N1965), .A(N1963), .B(N805), .CI(N704));
ADDFX1 inst_cellmath__203_0_I973 (.CO(N1968), .S(N1967), .A(N1938), .B(N732), .CI(N760));
ADDFX1 inst_cellmath__203_0_I974 (.CO(N1970), .S(N1969), .A(N1965), .B(N1940), .CI(N1942));
ADDFX1 inst_cellmath__203_0_I975 (.CO(inst_cellmath__203_0_out1[29]), .S(inst_cellmath__203_0_out0[28]), .A(N1944), .B(N1967), .CI(N1969));
ADDFX1 inst_cellmath__203_0_I976 (.CO(N1974), .S(N1973), .A(N1131), .B(N5720), .CI(N1221));
ADDFX1 inst_cellmath__203_0_I977 (.CO(N1976), .S(N1975), .A(N1251), .B(N1281), .CI(N1161));
ADDFX1 inst_cellmath__203_0_I978 (.CO(N1978), .S(N1977), .A(N1311), .B(N1191), .CI(N1948));
ADDFX1 inst_cellmath__203_0_I979 (.CO(N1980), .S(N1979), .A(N1954), .B(N1952), .CI(N1973));
ADDFX1 inst_cellmath__203_0_I980 (.CO(N1982), .S(N1981), .A(N1956), .B(N1975), .CI(N1977));
ADDFX1 inst_cellmath__203_0_I981 (.CO(N1984), .S(N1983), .A(N1958), .B(N1979), .CI(N1981));
ADDFX1 inst_cellmath__203_0_I982 (.CO(N1986), .S(N1985), .A(N1983), .B(N1960), .CI(N1962));
ADDFX1 inst_cellmath__203_0_I983 (.CO(N1988), .S(N1987), .A(N807), .B(N1985), .CI(N1964));
ADDFX1 inst_cellmath__203_0_I984 (.CO(N1990), .S(N1989), .A(N733), .B(N705), .CI(N761));
ADDFX1 inst_cellmath__203_0_I985 (.CO(N1992), .S(N1991), .A(N1966), .B(N1987), .CI(N1968));
ADDFX1 inst_cellmath__203_0_I986 (.CO(inst_cellmath__203_0_out1[30]), .S(inst_cellmath__203_0_out0[29]), .A(N1970), .B(N1989), .CI(N1991));
INVXL fap1_A_I1812 (.Y(N5518), .A(N5725));
ADDFX1 fap1_A_I1813 (.CO(N1996), .S(N1995), .A(N1282), .B(N1162), .CI(N5518));
ADDFX1 inst_cellmath__203_0_I988 (.CO(N2000), .S(N1999), .A(N1192), .B(N1252), .CI(N1222));
ADDFX1 inst_cellmath__203_0_I989 (.CO(N2002), .S(N2001), .A(N1974), .B(N1312), .CI(N1976));
ADDFX1 inst_cellmath__203_0_I990 (.CO(N2004), .S(N2003), .A(N1995), .B(N1978), .CI(N1999));
ADDFX1 inst_cellmath__203_0_I991 (.CO(N2006), .S(N2005), .A(N2001), .B(N1980), .CI(N1982));
ADDFX1 inst_cellmath__203_0_I992 (.CO(N2008), .S(N2007), .A(N1984), .B(N2003), .CI(N2005));
ADDFX1 inst_cellmath__203_0_I993 (.CO(N2010), .S(N2009), .A(N1986), .B(N2007), .CI(N5679));
ADDFX1 inst_cellmath__203_0_I994 (.CO(N2012), .S(N2011), .A(N2009), .B(N809), .CI(N734));
ADDFX1 inst_cellmath__203_0_I995 (.CO(N2014), .S(N2013), .A(N762), .B(N1988), .CI(N1990));
ADDFX1 inst_cellmath__203_0_I996 (.CO(inst_cellmath__203_0_out1[31]), .S(inst_cellmath__203_0_out0[30]), .A(N1992), .B(N2011), .CI(N2013));
ADDFX1 inst_cellmath__203_0_I997 (.CO(N2018), .S(N2017), .A(N1163), .B(N5725), .CI(N1253));
ADDFX1 inst_cellmath__203_0_I998 (.CO(N2020), .S(N2019), .A(N1283), .B(N1313), .CI(N1193));
ADDFX1 inst_cellmath__203_0_I999 (.CO(N2022), .S(N2021), .A(N1996), .B(N1223), .CI(N2000));
ADDFX1 inst_cellmath__203_0_I1000 (.CO(N2024), .S(N2023), .A(N2019), .B(N2017), .CI(N2002));
ADDFX1 inst_cellmath__203_0_I1001 (.CO(N2026), .S(N2025), .A(N2021), .B(N2004), .CI(N2023));
ADDFX1 inst_cellmath__203_0_I1002 (.CO(N2028), .S(N2027), .A(N2025), .B(N2006), .CI(N2008));
ADDFX1 inst_cellmath__203_0_I1003 (.CO(N2030), .S(N2029), .A(N811), .B(N2027), .CI(N2010));
ADDFX1 inst_cellmath__203_0_I1004 (.CO(N2032), .S(N2031), .A(N763), .B(N735), .CI(N2029));
ADDFX1 inst_cellmath__203_0_I1005 (.CO(inst_cellmath__203_0_out0[32]), .S(inst_cellmath__203_0_out0[31]), .A(N2031), .B(N2012), .CI(N2014));
INVXL fap1_A_I1814 (.Y(N5527), .A(N5730));
ADDFX1 fap1_A_I1815 (.CO(N2036), .S(N2035), .A(N1314), .B(N1194), .CI(N5527));
ADDFX1 inst_cellmath__203_0_I1007 (.CO(N2040), .S(N2039), .A(N1224), .B(N1284), .CI(N1254));
ADDFX1 inst_cellmath__203_0_I1008 (.CO(N2042), .S(N2041), .A(N2020), .B(N2018), .CI(N2035));
ADDFX1 inst_cellmath__203_0_I1009 (.CO(N2044), .S(N2043), .A(N2022), .B(N2039), .CI(N2024));
ADDFX1 inst_cellmath__203_0_I1010 (.CO(N2046), .S(N2045), .A(N2043), .B(N2041), .CI(N2026));
ADDFX1 inst_cellmath__203_0_I1011 (.CO(N2048), .S(N2047), .A(N2028), .B(N2045), .CI(N813));
ADDFX1 inst_cellmath__203_0_I1012 (.CO(N2050), .S(N2049), .A(N2030), .B(N5684), .CI(N2047));
ADDFX1 inst_cellmath__203_0_I1013 (.CO(inst_cellmath__203_0_out0[33]), .S(inst_cellmath__203_0_out1[32]), .A(N2049), .B(N764), .CI(N2032));
ADDFX1 inst_cellmath__203_0_I1014 (.CO(N2054), .S(N2053), .A(N1195), .B(N5730), .CI(N1285));
ADDFX1 inst_cellmath__203_0_I1015 (.CO(N2056), .S(N2055), .A(N1225), .B(N1315), .CI(N1255));
ADDFX1 inst_cellmath__203_0_I1016 (.CO(N2058), .S(N2057), .A(N2040), .B(N2036), .CI(N2053));
ADDFX1 inst_cellmath__203_0_I1017 (.CO(N2060), .S(N2059), .A(N2042), .B(N2055), .CI(N2057));
ADDFX1 inst_cellmath__203_0_I1018 (.CO(N2062), .S(N2061), .A(N2059), .B(N2044), .CI(N2046));
ADDFX1 inst_cellmath__203_0_I1019 (.CO(N2064), .S(N2063), .A(N815), .B(N2061), .CI(N2048));
ADDFX1 inst_cellmath__203_0_I1020 (.CO(inst_cellmath__203_0_out0[34]), .S(inst_cellmath__203_0_out1[33]), .A(N2063), .B(N765), .CI(N2050));
INVXL fap1_A_I1816 (.Y(N5536), .A(N5735));
ADDFX1 fap1_A_I1817 (.CO(N2068), .S(N2067), .A(N1316), .B(N1226), .CI(N5536));
ADDFX1 inst_cellmath__203_0_I1022 (.CO(N2072), .S(N2071), .A(N1286), .B(N1256), .CI(N2054));
ADDFX1 inst_cellmath__203_0_I1023 (.CO(N2074), .S(N2073), .A(N2067), .B(N2056), .CI(N2071));
ADDFX1 inst_cellmath__203_0_I1024 (.CO(N2076), .S(N2075), .A(N2060), .B(N2058), .CI(N2073));
ADDFX1 inst_cellmath__203_0_I1025 (.CO(N2078), .S(N2077), .A(N2062), .B(N2075), .CI(N817));
ADDFX1 inst_cellmath__203_0_I1026 (.CO(inst_cellmath__203_0_out0[35]), .S(inst_cellmath__203_0_out1[34]), .A(N2077), .B(N5689), .CI(N2064));
ADDFX1 inst_cellmath__203_0_I1027 (.CO(N2082), .S(N2081), .A(N1227), .B(N5735), .CI(N1317));
ADDFX1 inst_cellmath__203_0_I1028 (.CO(N2084), .S(N2083), .A(N1287), .B(N1257), .CI(N2068));
ADDFX1 inst_cellmath__203_0_I1029 (.CO(N2086), .S(N2085), .A(N2072), .B(N2081), .CI(N2083));
ADDFX1 inst_cellmath__203_0_I1030 (.CO(N2088), .S(N2087), .A(N2085), .B(N2074), .CI(N2076));
ADDFX1 inst_cellmath__203_0_I1031 (.CO(inst_cellmath__203_0_out0[36]), .S(inst_cellmath__203_0_out1[35]), .A(N819), .B(N2087), .CI(N2078));
INVXL fap1_A_I1818 (.Y(N5545), .A(N5740));
ADDFX1 fap1_A_I1819 (.CO(N2092), .S(N2091), .A(N1288), .B(N1258), .CI(N5545));
ADDFX1 inst_cellmath__203_0_I1033 (.CO(N2096), .S(N2095), .A(N2082), .B(N1318), .CI(N2091));
ADDFX1 inst_cellmath__203_0_I1034 (.CO(N2098), .S(N2097), .A(N2095), .B(N2084), .CI(N2086));
ADDFX1 inst_cellmath__203_0_I1035 (.CO(inst_cellmath__203_0_out0[37]), .S(inst_cellmath__203_0_out1[36]), .A(N2088), .B(N2097), .CI(N1366));
ADDFX1 inst_cellmath__203_0_I1036 (.CO(N2102), .S(N2101), .A(N1259), .B(N5740), .CI(N1289));
ADDFX1 inst_cellmath__203_0_I1037 (.CO(N2104), .S(N2103), .A(N2092), .B(N1319), .CI(N2101));
ADDFX1 inst_cellmath__203_0_I1038 (.CO(inst_cellmath__203_0_out0[38]), .S(inst_cellmath__203_0_out1[37]), .A(N2103), .B(N2096), .CI(N2098));
ADDFX1 inst_cellmath__203_0_I1039 (.CO(N2108), .S(N2107), .A(N1290), .B(N5745), .CI(N1320));
ADDFX1 inst_cellmath__203_0_I1040 (.CO(inst_cellmath__203_0_out0[39]), .S(inst_cellmath__203_0_out1[38]), .A(N2107), .B(N2102), .CI(N2104));
INVXL inst_cellmath__203_0_I1041 (.Y(N2111), .A(N2112));
ADDFX1 inst_cellmath__203_0_I1042 (.CO(inst_cellmath__203_0_out0[40]), .S(inst_cellmath__203_0_out1[39]), .A(N1321), .B(N2111), .CI(N2108));
ADDFX1 inst_cellmath__203_0_I1043 (.CO(inst_cellmath__203_0_out0[41]), .S(inst_cellmath__203_0_out1[40]), .A(N2112), .B(N5750), .CI(N1322));
INVXL inst_cellmath__203_0_I1044 (.Y(inst_cellmath__203_0_out1[41]), .A(inst_cellmath__203_0_out0[42]));
assign inst_cellmath__203_0_out0[0] = 1'B0;
assign inst_cellmath__203_0_out0[43] = 1'B0;
assign inst_cellmath__203_0_out0[44] = 1'B0;
assign inst_cellmath__203_0_out0[45] = 1'B0;
assign inst_cellmath__203_0_out0[46] = 1'B0;
assign inst_cellmath__203_0_out1[43] = 1'B1;
assign inst_cellmath__203_0_out1[44] = 1'B1;
assign inst_cellmath__203_0_out1[45] = 1'B1;
assign inst_cellmath__203_0_out1[46] = 1'B1;
endmodule

module cynw_cm_float_cos_inst_cellmath__201_0_bdw1114505291_bdw (
	inst_cellmath__201_0_out0,
	inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1,
	inst_cellmath__201_0_in2
	); /* architecture "gate_level" */ 
output [49:0] inst_cellmath__201_0_out0;
input [46:0] inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1;
input [72:43] inst_cellmath__201_0_in2;
wire [46:0] inst_cellmath__203__W1;
wire N989,N991,N992,N993,N994,N995,N996 
	,N997,N998,N999,N1000,N1001,N1002,N1003,N1004 
	,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012 
	,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020 
	,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028 
	,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036 
	,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044 
	,N1045,N1046,N1047,N1048,N1049,N1053,N1054,N1055 
	,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063 
	,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071 
	,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079 
	,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087 
	,N1088,N1089,N1090,N1091,N1094,N1102,N1110,N1122 
	,N1134,N1150,N1166,N1186,N1206,N1230,N1254,N1282 
	,N1318,N1320,N1324,N1325,N1328,N1329,N1382,N1449 
	,N1452,N1455,N1458,N1461,N1464,N1467,N1470,N1473 
	,N1476,N1479,N1482,N1485,N1488,N1491,N1494,N1497 
	,N1500,N1503,N1524,N1526,N1527,N1528,N1529,N1530 
	,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538 
	,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546 
	,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554 
	,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562 
	,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570 
	,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578 
	,N1579,N1580,N1581,N1585,N1587,N1588,N1589,N1590 
	,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598 
	,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606 
	,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614 
	,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622 
	,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630 
	,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638 
	,N1639,N1640,N1643,N1648,N1650,N1652,N1653,N1654 
	,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662 
	,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670 
	,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678 
	,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686 
	,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694 
	,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702 
	,N1703,N1712,N1714,N1716,N1718,N1720,N1721,N1722 
	,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730 
	,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738 
	,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746 
	,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754 
	,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762 
	,N1763,N1780,N1782,N1784,N1786,N1788,N1790,N1796 
	,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804 
	,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812 
	,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820 
	,N1821,N1822,N1823,N1856,N1858,N1860,N1862,N1864 
	,N1866,N1868,N1870,N1872,N1874,N1876,N1878,N1880 
	,N1889,N1892,N1895,N1898,N1901,N1904,N1907,N1910 
	,N1913,N1916,N1919,N1922,N1925,N1928,N1931,N1934 
	,N1937,N1940,N1943,N1946,N1949,N1952,N1955,N1958 
	,N1961,N1964,N1967,N1970,N2234,N2235,N2241,N2242 
	,N2252,N2253,N2267,N2268,N2286,N2287,N2309,N2310 
	,N2329,N2349,N2358,N2359,N2392,N2393,N2394,N2440 
	,N2441,N2493,N2502,N2504,N2510;
INVXL inst_cellmath__201_0_I102 (.Y(inst_cellmath__203__W1[46]), .A(inst_cellmath__201_0_in0[46]));
INVXL inst_cellmath__201_0_I243 (.Y(N989), .A(inst_cellmath__201_0_in1[46]));
ADDHX1 inst_cellmath__201_0_I245 (.CO(N992), .S(N991), .A(inst_cellmath__201_0_in2[43]), .B(inst_cellmath__201_0_in1[18]));
ADDFX1 inst_cellmath__201_0_I246 (.CO(N994), .S(N993), .A(inst_cellmath__201_0_in1[19]), .B(inst_cellmath__201_0_in2[44]), .CI(inst_cellmath__201_0_in0[19]));
ADDFX1 inst_cellmath__201_0_I247 (.CO(N996), .S(N995), .A(inst_cellmath__201_0_in1[20]), .B(inst_cellmath__201_0_in2[45]), .CI(inst_cellmath__201_0_in0[20]));
ADDFX1 inst_cellmath__201_0_I248 (.CO(N998), .S(N997), .A(inst_cellmath__201_0_in1[21]), .B(inst_cellmath__201_0_in2[46]), .CI(inst_cellmath__201_0_in0[21]));
ADDFX1 inst_cellmath__201_0_I249 (.CO(N1000), .S(N999), .A(inst_cellmath__201_0_in1[22]), .B(inst_cellmath__201_0_in2[47]), .CI(inst_cellmath__201_0_in0[22]));
ADDFX1 inst_cellmath__201_0_I250 (.CO(N1002), .S(N1001), .A(inst_cellmath__201_0_in1[23]), .B(inst_cellmath__201_0_in2[48]), .CI(inst_cellmath__201_0_in0[23]));
ADDFX1 inst_cellmath__201_0_I251 (.CO(N1004), .S(N1003), .A(inst_cellmath__201_0_in1[24]), .B(inst_cellmath__201_0_in2[49]), .CI(inst_cellmath__201_0_in0[24]));
ADDFX1 inst_cellmath__201_0_I252 (.CO(N1006), .S(N1005), .A(inst_cellmath__201_0_in1[25]), .B(inst_cellmath__201_0_in2[50]), .CI(inst_cellmath__201_0_in0[25]));
ADDFX1 inst_cellmath__201_0_I253 (.CO(N1008), .S(N1007), .A(inst_cellmath__201_0_in1[26]), .B(inst_cellmath__201_0_in2[51]), .CI(inst_cellmath__201_0_in0[26]));
ADDFX1 inst_cellmath__201_0_I254 (.CO(N1010), .S(N1009), .A(inst_cellmath__201_0_in1[27]), .B(inst_cellmath__201_0_in2[52]), .CI(inst_cellmath__201_0_in0[27]));
ADDFX1 inst_cellmath__201_0_I255 (.CO(N1012), .S(N1011), .A(inst_cellmath__201_0_in1[28]), .B(inst_cellmath__201_0_in2[53]), .CI(inst_cellmath__201_0_in0[28]));
ADDFX1 inst_cellmath__201_0_I256 (.CO(N1014), .S(N1013), .A(inst_cellmath__201_0_in1[29]), .B(inst_cellmath__201_0_in2[54]), .CI(inst_cellmath__201_0_in0[29]));
ADDFX1 inst_cellmath__201_0_I257 (.CO(N1016), .S(N1015), .A(inst_cellmath__201_0_in1[30]), .B(inst_cellmath__201_0_in2[55]), .CI(inst_cellmath__201_0_in0[30]));
ADDFX1 inst_cellmath__201_0_I258 (.CO(N1018), .S(N1017), .A(inst_cellmath__201_0_in1[31]), .B(inst_cellmath__201_0_in2[56]), .CI(inst_cellmath__201_0_in0[31]));
ADDFX1 inst_cellmath__201_0_I259 (.CO(N1020), .S(N1019), .A(inst_cellmath__201_0_in1[32]), .B(inst_cellmath__201_0_in2[57]), .CI(inst_cellmath__201_0_in0[32]));
ADDFX1 inst_cellmath__201_0_I260 (.CO(N1022), .S(N1021), .A(inst_cellmath__201_0_in0[33]), .B(inst_cellmath__201_0_in2[58]), .CI(inst_cellmath__201_0_in1[33]));
ADDFX1 inst_cellmath__201_0_I261 (.CO(N1024), .S(N1023), .A(inst_cellmath__201_0_in1[34]), .B(inst_cellmath__201_0_in2[59]), .CI(inst_cellmath__201_0_in0[34]));
ADDFX1 inst_cellmath__201_0_I262 (.CO(N1026), .S(N1025), .A(inst_cellmath__201_0_in0[35]), .B(inst_cellmath__201_0_in2[60]), .CI(inst_cellmath__201_0_in1[35]));
ADDFX1 inst_cellmath__201_0_I263 (.CO(N1028), .S(N1027), .A(inst_cellmath__201_0_in1[36]), .B(inst_cellmath__201_0_in2[61]), .CI(inst_cellmath__201_0_in0[36]));
ADDFX1 inst_cellmath__201_0_I264 (.CO(N1030), .S(N1029), .A(inst_cellmath__201_0_in1[37]), .B(inst_cellmath__201_0_in2[62]), .CI(inst_cellmath__201_0_in0[37]));
ADDFX1 inst_cellmath__201_0_I265 (.CO(N1032), .S(N1031), .A(inst_cellmath__201_0_in1[38]), .B(inst_cellmath__201_0_in2[63]), .CI(inst_cellmath__201_0_in0[38]));
ADDFX1 inst_cellmath__201_0_I266 (.CO(N1034), .S(N1033), .A(inst_cellmath__201_0_in1[39]), .B(inst_cellmath__201_0_in2[64]), .CI(inst_cellmath__201_0_in0[39]));
ADDFX1 inst_cellmath__201_0_I267 (.CO(N1036), .S(N1035), .A(inst_cellmath__201_0_in1[40]), .B(inst_cellmath__201_0_in2[65]), .CI(inst_cellmath__201_0_in0[40]));
ADDFX1 inst_cellmath__201_0_I268 (.CO(N1038), .S(N1037), .A(inst_cellmath__201_0_in2[66]), .B(inst_cellmath__201_0_in1[41]), .CI(inst_cellmath__201_0_in0[41]));
ADDFX1 inst_cellmath__201_0_I269 (.CO(N1040), .S(N1039), .A(inst_cellmath__201_0_in0[42]), .B(inst_cellmath__201_0_in1[42]), .CI(inst_cellmath__201_0_in2[67]));
ADDFX1 inst_cellmath__201_0_I270 (.CO(N1042), .S(N1041), .A(inst_cellmath__201_0_in0[43]), .B(inst_cellmath__201_0_in1[43]), .CI(inst_cellmath__201_0_in2[68]));
ADDFX1 inst_cellmath__201_0_I271 (.CO(N1044), .S(N1043), .A(inst_cellmath__201_0_in0[44]), .B(inst_cellmath__201_0_in1[44]), .CI(inst_cellmath__201_0_in2[69]));
ADDFX1 inst_cellmath__201_0_I272 (.CO(N1046), .S(N1045), .A(inst_cellmath__201_0_in0[45]), .B(inst_cellmath__201_0_in1[45]), .CI(inst_cellmath__201_0_in2[70]));
ADDFX1 inst_cellmath__201_0_I273 (.CO(N1048), .S(N1047), .A(inst_cellmath__203__W1[46]), .B(N989), .CI(inst_cellmath__201_0_in2[71]));
INVXL inst_cellmath__201_0_I274 (.Y(N1049), .A(inst_cellmath__201_0_in2[72]));
NAND2XL inst_cellmath__201_0_I275 (.Y(N1053), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
NOR2XL inst_cellmath__201_0_I276 (.Y(N1054), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NAND2XL inst_cellmath__201_0_I277 (.Y(N1055), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NOR2XL inst_cellmath__201_0_I278 (.Y(N1056), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NAND2XL inst_cellmath__201_0_I279 (.Y(N1057), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NOR2XL inst_cellmath__201_0_I280 (.Y(N1058), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NAND2XL inst_cellmath__201_0_I281 (.Y(N1059), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NOR2XL inst_cellmath__201_0_I282 (.Y(N1060), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NAND2XL inst_cellmath__201_0_I283 (.Y(N1061), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NOR2XL inst_cellmath__201_0_I284 (.Y(N1062), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NAND2XL inst_cellmath__201_0_I285 (.Y(N1063), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NOR2XL inst_cellmath__201_0_I286 (.Y(N1064), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NAND2XL inst_cellmath__201_0_I287 (.Y(N1065), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NOR2XL inst_cellmath__201_0_I288 (.Y(N1066), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NAND2XL inst_cellmath__201_0_I289 (.Y(N1067), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NOR2XL inst_cellmath__201_0_I290 (.Y(N1068), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NAND2XL inst_cellmath__201_0_I291 (.Y(N1069), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NOR2XL inst_cellmath__201_0_I292 (.Y(N1070), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NAND2XL inst_cellmath__201_0_I293 (.Y(N1071), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NOR2XL inst_cellmath__201_0_I294 (.Y(N1072), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NAND2XL inst_cellmath__201_0_I295 (.Y(N1073), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NOR2XL inst_cellmath__201_0_I296 (.Y(N1074), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NAND2XL inst_cellmath__201_0_I297 (.Y(N1075), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NOR2XL inst_cellmath__201_0_I298 (.Y(N1076), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NAND2XL inst_cellmath__201_0_I299 (.Y(N1077), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NOR2XL inst_cellmath__201_0_I300 (.Y(N1078), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NAND2XL inst_cellmath__201_0_I301 (.Y(N1079), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NOR2XL inst_cellmath__201_0_I302 (.Y(N1080), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NAND2XL inst_cellmath__201_0_I303 (.Y(N1081), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NOR2XL inst_cellmath__201_0_I304 (.Y(N1082), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NAND2XL inst_cellmath__201_0_I305 (.Y(N1083), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NOR2XL inst_cellmath__201_0_I306 (.Y(N1084), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
NAND2XL inst_cellmath__201_0_I307 (.Y(N1085), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
NOR2XL inst_cellmath__201_0_I308 (.Y(N1086), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NAND2XL inst_cellmath__201_0_I309 (.Y(N1087), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NOR2XL inst_cellmath__201_0_I310 (.Y(N1088), .A(inst_cellmath__201_0_in0[18]), .B(N991));
NAND2XL inst_cellmath__201_0_I311 (.Y(N1089), .A(inst_cellmath__201_0_in0[18]), .B(N991));
NOR2XL inst_cellmath__201_0_I312 (.Y(N1090), .A(N992), .B(N993));
NAND2XL inst_cellmath__201_0_I313 (.Y(N1091), .A(N992), .B(N993));
AOI21XL inst_cellmath__201_0_I316 (.Y(N1094), .A0(N1055), .A1(N1053), .B0(N1054));
INVXL inst_cellmath__201_0_I1343 (.Y(N2234), .A(N1056));
INVXL inst_cellmath__201_0_I1344 (.Y(N2235), .A(N1057));
OAI21XL inst_cellmath__201_0_I324 (.Y(N1102), .A0(N2235), .A1(N1094), .B0(N2234));
AOI21XL inst_cellmath__201_0_I332 (.Y(N1110), .A0(N1059), .A1(N1102), .B0(N1058));
INVXL inst_cellmath__201_0_I1350 (.Y(N2241), .A(N1060));
INVXL inst_cellmath__201_0_I1351 (.Y(N2242), .A(N1061));
OAI21XL inst_cellmath__201_0_I344 (.Y(N1122), .A0(N2242), .A1(N1110), .B0(N2241));
AOI21XL inst_cellmath__201_0_I356 (.Y(N1134), .A0(N1063), .A1(N1122), .B0(N1062));
INVXL inst_cellmath__201_0_I1361 (.Y(N2252), .A(N1064));
INVXL inst_cellmath__201_0_I1362 (.Y(N2253), .A(N1065));
OAI21XL inst_cellmath__201_0_I372 (.Y(N1150), .A0(N2253), .A1(N1134), .B0(N2252));
AOI21XL inst_cellmath__201_0_I388 (.Y(N1166), .A0(N1067), .A1(N1150), .B0(N1066));
INVXL inst_cellmath__201_0_I1376 (.Y(N2267), .A(N1068));
INVXL inst_cellmath__201_0_I1377 (.Y(N2268), .A(N1069));
OAI21XL inst_cellmath__201_0_I408 (.Y(N1186), .A0(N2268), .A1(N1166), .B0(N2267));
AOI21XL inst_cellmath__201_0_I428 (.Y(N1206), .A0(N1071), .A1(N1186), .B0(N1070));
INVXL inst_cellmath__201_0_I1395 (.Y(N2286), .A(N1072));
INVXL inst_cellmath__201_0_I1396 (.Y(N2287), .A(N1073));
OAI21XL inst_cellmath__201_0_I452 (.Y(N1230), .A0(N2287), .A1(N1206), .B0(N2286));
AOI21XL inst_cellmath__201_0_I476 (.Y(N1254), .A0(N1075), .A1(N1230), .B0(N1074));
INVXL inst_cellmath__201_0_I1418 (.Y(N2309), .A(N1076));
INVXL inst_cellmath__201_0_I1419 (.Y(N2310), .A(N1077));
OAI21XL inst_cellmath__201_0_I504 (.Y(N1282), .A0(N2310), .A1(N1254), .B0(N2309));
AO21XL inst_cellmath__201_0_I1566 (.Y(N2329), .A0(N1081), .A1(N1078), .B0(N1080));
AOI21XL inst_cellmath__201_0_I540 (.Y(N1318), .A0(N1079), .A1(N1282), .B0(N1078));
AOI31X1 inst_cellmath__201_0_I2623 (.Y(N1320), .A0(N1081), .A1(N1079), .A2(N1282), .B0(N2329));
AOI21XL inst_cellmath__201_0_I546 (.Y(N1324), .A0(N1085), .A1(N1082), .B0(N1084));
NAND2XL inst_cellmath__201_0_I547 (.Y(N1325), .A(N1085), .B(N1083));
INVXL inst_cellmath__201_0_I1458 (.Y(N2349), .A(N1087));
AOI21XL inst_cellmath__201_0_I550 (.Y(N1328), .A0(N1089), .A1(N1086), .B0(N1088));
NAND2XL inst_cellmath__201_0_I551 (.Y(N1329), .A(N1089), .B(N1087));
NOR2XL andori2bb1_A_I1638 (.Y(N2493), .A(N2349), .B(N1324));
NOR2XL andori2bb1_A_I1639 (.Y(N2358), .A(N2493), .B(N1086));
OR2XL inst_cellmath__201_0_I1570 (.Y(N2359), .A(N2349), .B(N1325));
OAI21XL orandi31_A_I2624 (.Y(N2504), .A0(N1329), .A1(N1324), .B0(N1328));
NOR3XL orandi31_A_I1641 (.Y(N2502), .A(N1329), .B(N1325), .C(N1320));
OR2XL orandi31_A_I1642 (.Y(N1382), .A(N2502), .B(N2504));
NOR2BX1 andori2bb1_A_I2625 (.Y(N2510), .AN(N1083), .B(N1320));
NOR2XL andori2bb1_A_I1644 (.Y(N2392), .A(N2510), .B(N1082));
OA21X1 inst_cellmath__201_0_I1576 (.Y(N2393), .A0(N1325), .A1(N1320), .B0(N1324));
OA21X1 inst_cellmath__201_0_I1577 (.Y(N2394), .A0(N2359), .A1(N1320), .B0(N2358));
NAND2BXL inst_cellmath__201_0_I671 (.Y(N1449), .AN(N1054), .B(N1055));
NAND2BXL inst_cellmath__201_0_I674 (.Y(N1452), .AN(N1056), .B(N1057));
NAND2BXL inst_cellmath__201_0_I677 (.Y(N1455), .AN(N1058), .B(N1059));
NAND2BXL inst_cellmath__201_0_I680 (.Y(N1458), .AN(N1060), .B(N1061));
NAND2BXL inst_cellmath__201_0_I683 (.Y(N1461), .AN(N1062), .B(N1063));
NAND2BXL inst_cellmath__201_0_I686 (.Y(N1464), .AN(N1064), .B(N1065));
NAND2BXL inst_cellmath__201_0_I689 (.Y(N1467), .AN(N1066), .B(N1067));
NAND2BXL inst_cellmath__201_0_I692 (.Y(N1470), .AN(N1068), .B(N1069));
NAND2BXL inst_cellmath__201_0_I695 (.Y(N1473), .AN(N1070), .B(N1071));
NAND2BXL inst_cellmath__201_0_I698 (.Y(N1476), .AN(N1072), .B(N1073));
NAND2BXL inst_cellmath__201_0_I701 (.Y(N1479), .AN(N1074), .B(N1075));
NAND2BXL inst_cellmath__201_0_I704 (.Y(N1482), .AN(N1076), .B(N1077));
NAND2BXL inst_cellmath__201_0_I707 (.Y(N1485), .AN(N1078), .B(N1079));
NAND2BXL inst_cellmath__201_0_I710 (.Y(N1488), .AN(N1080), .B(N1081));
NAND2BXL inst_cellmath__201_0_I713 (.Y(N1491), .AN(N1082), .B(N1083));
NAND2BXL inst_cellmath__201_0_I716 (.Y(N1494), .AN(N1084), .B(N1085));
NAND2BXL inst_cellmath__201_0_I719 (.Y(N1497), .AN(N1086), .B(N1087));
NAND2BXL inst_cellmath__201_0_I722 (.Y(N1500), .AN(N1088), .B(N1089));
NAND2BXL inst_cellmath__201_0_I725 (.Y(N1503), .AN(N1090), .B(N1091));
XOR2XL inst_cellmath__201_0_I2626 (.Y(inst_cellmath__201_0_out0[0]), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
XOR2XL inst_cellmath__201_0_I2627 (.Y(inst_cellmath__201_0_out0[1]), .A(N1053), .B(N1449));
XNOR2X1 inst_cellmath__201_0_I1579 (.Y(inst_cellmath__201_0_out0[2]), .A(N1094), .B(N1452));
XOR2XL inst_cellmath__201_0_I1612 (.Y(inst_cellmath__201_0_out0[3]), .A(N1102), .B(N1455));
XNOR2X1 inst_cellmath__201_0_I1581 (.Y(inst_cellmath__201_0_out0[4]), .A(N1110), .B(N1458));
XOR2XL inst_cellmath__201_0_I1582 (.Y(inst_cellmath__201_0_out0[5]), .A(N1122), .B(N1461));
XNOR2X1 inst_cellmath__201_0_I732 (.Y(inst_cellmath__201_0_out0[6]), .A(N1134), .B(N1464));
XOR2XL inst_cellmath__201_0_I1583 (.Y(inst_cellmath__201_0_out0[7]), .A(N1150), .B(N1467));
XNOR2X1 inst_cellmath__201_0_I734 (.Y(inst_cellmath__201_0_out0[8]), .A(N1166), .B(N1470));
XOR2XL inst_cellmath__201_0_I1584 (.Y(inst_cellmath__201_0_out0[9]), .A(N1186), .B(N1473));
XNOR2X1 inst_cellmath__201_0_I736 (.Y(inst_cellmath__201_0_out0[10]), .A(N1206), .B(N1476));
XOR2XL inst_cellmath__201_0_I1585 (.Y(inst_cellmath__201_0_out0[11]), .A(N1230), .B(N1479));
XNOR2X1 inst_cellmath__201_0_I738 (.Y(inst_cellmath__201_0_out0[12]), .A(N1254), .B(N1482));
XOR2XL inst_cellmath__201_0_I1586 (.Y(inst_cellmath__201_0_out0[13]), .A(N1282), .B(N1485));
XNOR2X1 inst_cellmath__201_0_I740 (.Y(inst_cellmath__201_0_out0[14]), .A(N1318), .B(N1488));
XNOR2X1 inst_cellmath__201_0_I741 (.Y(inst_cellmath__201_0_out0[15]), .A(N1320), .B(N1491));
XNOR2X1 inst_cellmath__201_0_I742 (.Y(inst_cellmath__201_0_out0[16]), .A(N2392), .B(N1494));
XNOR2X1 inst_cellmath__201_0_I743 (.Y(inst_cellmath__201_0_out0[17]), .A(N2393), .B(N1497));
XNOR2X1 inst_cellmath__201_0_I744 (.Y(inst_cellmath__201_0_out0[18]), .A(N2394), .B(N1500));
XOR2XL inst_cellmath__201_0_I1587 (.Y(inst_cellmath__201_0_out0[19]), .A(N1382), .B(N1503));
AO21XL inst_cellmath__201_0_I1613 (.Y(N1524), .A0(N1091), .A1(N1382), .B0(N1090));
NOR2XL inst_cellmath__201_0_I747 (.Y(N1526), .A(N994), .B(N995));
NAND2XL inst_cellmath__201_0_I748 (.Y(N1527), .A(N994), .B(N995));
NOR2XL inst_cellmath__201_0_I749 (.Y(N1528), .A(N996), .B(N997));
NAND2XL inst_cellmath__201_0_I750 (.Y(N1529), .A(N996), .B(N997));
NOR2XL inst_cellmath__201_0_I751 (.Y(N1530), .A(N998), .B(N999));
NAND2XL inst_cellmath__201_0_I752 (.Y(N1531), .A(N998), .B(N999));
NOR2XL inst_cellmath__201_0_I753 (.Y(N1532), .A(N1000), .B(N1001));
NAND2XL inst_cellmath__201_0_I754 (.Y(N1533), .A(N1000), .B(N1001));
NOR2XL inst_cellmath__201_0_I755 (.Y(N1534), .A(N1002), .B(N1003));
NAND2XL inst_cellmath__201_0_I756 (.Y(N1535), .A(N1002), .B(N1003));
NOR2XL inst_cellmath__201_0_I757 (.Y(N1536), .A(N1004), .B(N1005));
NAND2XL inst_cellmath__201_0_I758 (.Y(N1537), .A(N1004), .B(N1005));
NOR2XL inst_cellmath__201_0_I759 (.Y(N1538), .A(N1006), .B(N1007));
NAND2XL inst_cellmath__201_0_I760 (.Y(N1539), .A(N1006), .B(N1007));
NOR2XL inst_cellmath__201_0_I761 (.Y(N1540), .A(N1008), .B(N1009));
NAND2XL inst_cellmath__201_0_I762 (.Y(N1541), .A(N1008), .B(N1009));
NOR2XL inst_cellmath__201_0_I763 (.Y(N1542), .A(N1010), .B(N1011));
NAND2XL inst_cellmath__201_0_I764 (.Y(N1543), .A(N1010), .B(N1011));
NOR2XL inst_cellmath__201_0_I765 (.Y(N1544), .A(N1012), .B(N1013));
NAND2XL inst_cellmath__201_0_I766 (.Y(N1545), .A(N1012), .B(N1013));
NOR2XL inst_cellmath__201_0_I767 (.Y(N1546), .A(N1014), .B(N1015));
NAND2XL inst_cellmath__201_0_I768 (.Y(N1547), .A(N1014), .B(N1015));
NOR2XL inst_cellmath__201_0_I769 (.Y(N1548), .A(N1016), .B(N1017));
NAND2XL inst_cellmath__201_0_I770 (.Y(N1549), .A(N1016), .B(N1017));
NOR2XL inst_cellmath__201_0_I771 (.Y(N1550), .A(N1018), .B(N1019));
NAND2XL inst_cellmath__201_0_I772 (.Y(N1551), .A(N1018), .B(N1019));
NOR2XL inst_cellmath__201_0_I773 (.Y(N1552), .A(N1020), .B(N1021));
NAND2XL inst_cellmath__201_0_I774 (.Y(N1553), .A(N1020), .B(N1021));
NOR2XL inst_cellmath__201_0_I775 (.Y(N1554), .A(N1022), .B(N1023));
NAND2XL inst_cellmath__201_0_I776 (.Y(N1555), .A(N1022), .B(N1023));
NOR2XL inst_cellmath__201_0_I777 (.Y(N1556), .A(N1024), .B(N1025));
NAND2XL inst_cellmath__201_0_I778 (.Y(N1557), .A(N1024), .B(N1025));
NOR2XL inst_cellmath__201_0_I779 (.Y(N1558), .A(N1027), .B(N1026));
NAND2XL inst_cellmath__201_0_I780 (.Y(N1559), .A(N1027), .B(N1026));
NOR2XL inst_cellmath__201_0_I781 (.Y(N1560), .A(N1029), .B(N1028));
NAND2XL inst_cellmath__201_0_I782 (.Y(N1561), .A(N1029), .B(N1028));
NOR2XL inst_cellmath__201_0_I783 (.Y(N1562), .A(N1031), .B(N1030));
NAND2XL inst_cellmath__201_0_I784 (.Y(N1563), .A(N1031), .B(N1030));
NOR2XL inst_cellmath__201_0_I785 (.Y(N1564), .A(N1033), .B(N1032));
NAND2XL inst_cellmath__201_0_I786 (.Y(N1565), .A(N1033), .B(N1032));
NOR2XL inst_cellmath__201_0_I787 (.Y(N1566), .A(N1035), .B(N1034));
NAND2XL inst_cellmath__201_0_I788 (.Y(N1567), .A(N1035), .B(N1034));
NOR2XL inst_cellmath__201_0_I789 (.Y(N1568), .A(N1037), .B(N1036));
NAND2XL inst_cellmath__201_0_I790 (.Y(N1569), .A(N1037), .B(N1036));
NOR2XL inst_cellmath__201_0_I791 (.Y(N1570), .A(N1039), .B(N1038));
NAND2XL inst_cellmath__201_0_I792 (.Y(N1571), .A(N1039), .B(N1038));
NOR2XL inst_cellmath__201_0_I793 (.Y(N1572), .A(N1040), .B(N1041));
NAND2XL inst_cellmath__201_0_I794 (.Y(N1573), .A(N1040), .B(N1041));
NOR2XL inst_cellmath__201_0_I795 (.Y(N1574), .A(N1042), .B(N1043));
NAND2XL inst_cellmath__201_0_I796 (.Y(N1575), .A(N1042), .B(N1043));
NOR2XL inst_cellmath__201_0_I797 (.Y(N1576), .A(N1044), .B(N1045));
NAND2XL inst_cellmath__201_0_I798 (.Y(N1577), .A(N1044), .B(N1045));
NOR2XL inst_cellmath__201_0_I799 (.Y(N1578), .A(N1047), .B(N1046));
NAND2XL inst_cellmath__201_0_I800 (.Y(N1579), .A(N1047), .B(N1046));
NOR2XL inst_cellmath__201_0_I801 (.Y(N1580), .A(N1049), .B(N1048));
NAND2XL inst_cellmath__201_0_I802 (.Y(N1581), .A(N1049), .B(N1048));
AO21XL inst_cellmath__201_0_I806 (.Y(N1585), .A0(N1527), .A1(N1524), .B0(N1526));
AO21XL inst_cellmath__201_0_I808 (.Y(N1587), .A0(N1529), .A1(N1526), .B0(N1528));
AND2XL inst_cellmath__201_0_I809 (.Y(N1588), .A(N1529), .B(N1527));
AO21XL inst_cellmath__201_0_I810 (.Y(N1589), .A0(N1531), .A1(N1528), .B0(N1530));
AND2XL inst_cellmath__201_0_I811 (.Y(N1590), .A(N1531), .B(N1529));
AO21XL inst_cellmath__201_0_I812 (.Y(N1591), .A0(N1533), .A1(N1530), .B0(N1532));
AND2XL inst_cellmath__201_0_I813 (.Y(N1592), .A(N1533), .B(N1531));
AO21XL inst_cellmath__201_0_I814 (.Y(N1593), .A0(N1535), .A1(N1532), .B0(N1534));
AND2XL inst_cellmath__201_0_I815 (.Y(N1594), .A(N1535), .B(N1533));
AO21XL inst_cellmath__201_0_I816 (.Y(N1595), .A0(N1537), .A1(N1534), .B0(N1536));
AND2XL inst_cellmath__201_0_I817 (.Y(N1596), .A(N1537), .B(N1535));
AO21XL inst_cellmath__201_0_I818 (.Y(N1597), .A0(N1539), .A1(N1536), .B0(N1538));
AND2XL inst_cellmath__201_0_I819 (.Y(N1598), .A(N1539), .B(N1537));
AO21XL inst_cellmath__201_0_I820 (.Y(N1599), .A0(N1541), .A1(N1538), .B0(N1540));
AND2XL inst_cellmath__201_0_I821 (.Y(N1600), .A(N1541), .B(N1539));
AO21XL inst_cellmath__201_0_I822 (.Y(N1601), .A0(N1543), .A1(N1540), .B0(N1542));
AND2XL inst_cellmath__201_0_I823 (.Y(N1602), .A(N1543), .B(N1541));
AO21XL inst_cellmath__201_0_I824 (.Y(N1603), .A0(N1545), .A1(N1542), .B0(N1544));
AND2XL inst_cellmath__201_0_I825 (.Y(N1604), .A(N1545), .B(N1543));
AO21XL inst_cellmath__201_0_I826 (.Y(N1605), .A0(N1547), .A1(N1544), .B0(N1546));
AND2XL inst_cellmath__201_0_I827 (.Y(N1606), .A(N1547), .B(N1545));
AO21XL inst_cellmath__201_0_I828 (.Y(N1607), .A0(N1549), .A1(N1546), .B0(N1548));
AND2XL inst_cellmath__201_0_I829 (.Y(N1608), .A(N1549), .B(N1547));
AO21XL inst_cellmath__201_0_I830 (.Y(N1609), .A0(N1551), .A1(N1548), .B0(N1550));
AND2XL inst_cellmath__201_0_I831 (.Y(N1610), .A(N1551), .B(N1549));
AO21XL inst_cellmath__201_0_I832 (.Y(N1611), .A0(N1553), .A1(N1550), .B0(N1552));
AND2XL inst_cellmath__201_0_I833 (.Y(N1612), .A(N1553), .B(N1551));
AO21XL inst_cellmath__201_0_I834 (.Y(N1613), .A0(N1555), .A1(N1552), .B0(N1554));
AND2XL inst_cellmath__201_0_I835 (.Y(N1614), .A(N1555), .B(N1553));
AO21XL inst_cellmath__201_0_I836 (.Y(N1615), .A0(N1557), .A1(N1554), .B0(N1556));
AND2XL inst_cellmath__201_0_I837 (.Y(N1616), .A(N1557), .B(N1555));
AO21XL inst_cellmath__201_0_I838 (.Y(N1617), .A0(N1559), .A1(N1556), .B0(N1558));
AND2XL inst_cellmath__201_0_I839 (.Y(N1618), .A(N1559), .B(N1557));
AO21XL inst_cellmath__201_0_I840 (.Y(N1619), .A0(N1561), .A1(N1558), .B0(N1560));
AND2XL inst_cellmath__201_0_I841 (.Y(N1620), .A(N1561), .B(N1559));
AO21XL inst_cellmath__201_0_I842 (.Y(N1621), .A0(N1563), .A1(N1560), .B0(N1562));
AND2XL inst_cellmath__201_0_I843 (.Y(N1622), .A(N1563), .B(N1561));
AO21XL inst_cellmath__201_0_I844 (.Y(N1623), .A0(N1565), .A1(N1562), .B0(N1564));
AND2XL inst_cellmath__201_0_I845 (.Y(N1624), .A(N1565), .B(N1563));
AO21XL inst_cellmath__201_0_I846 (.Y(N1625), .A0(N1567), .A1(N1564), .B0(N1566));
AND2XL inst_cellmath__201_0_I847 (.Y(N1626), .A(N1567), .B(N1565));
AO21XL inst_cellmath__201_0_I848 (.Y(N1627), .A0(N1569), .A1(N1566), .B0(N1568));
AND2XL inst_cellmath__201_0_I849 (.Y(N1628), .A(N1569), .B(N1567));
AO21XL inst_cellmath__201_0_I850 (.Y(N1629), .A0(N1571), .A1(N1568), .B0(N1570));
AND2XL inst_cellmath__201_0_I851 (.Y(N1630), .A(N1571), .B(N1569));
AO21XL inst_cellmath__201_0_I852 (.Y(N1631), .A0(N1573), .A1(N1570), .B0(N1572));
AND2XL inst_cellmath__201_0_I853 (.Y(N1632), .A(N1573), .B(N1571));
AO21XL inst_cellmath__201_0_I854 (.Y(N1633), .A0(N1575), .A1(N1572), .B0(N1574));
AND2XL inst_cellmath__201_0_I855 (.Y(N1634), .A(N1575), .B(N1573));
AO21XL inst_cellmath__201_0_I856 (.Y(N1635), .A0(N1577), .A1(N1574), .B0(N1576));
AND2XL inst_cellmath__201_0_I857 (.Y(N1636), .A(N1577), .B(N1575));
AO21XL inst_cellmath__201_0_I858 (.Y(N1637), .A0(N1579), .A1(N1576), .B0(N1578));
AND2XL inst_cellmath__201_0_I859 (.Y(N1638), .A(N1579), .B(N1577));
AO21XL inst_cellmath__201_0_I860 (.Y(N1639), .A0(N1581), .A1(N1578), .B0(N1580));
AND2XL inst_cellmath__201_0_I861 (.Y(N1640), .A(N1581), .B(N1579));
AND2XL inst_cellmath__201_0_I863 (.Y(N1643), .A(N1049), .B(N1581));
AO21XL inst_cellmath__201_0_I868 (.Y(N1648), .A0(N1588), .A1(N1524), .B0(N1587));
AO21XL inst_cellmath__201_0_I870 (.Y(N1650), .A0(N1590), .A1(N1585), .B0(N1589));
AO21XL inst_cellmath__201_0_I872 (.Y(N1652), .A0(N1592), .A1(N1587), .B0(N1591));
AND2XL inst_cellmath__201_0_I873 (.Y(N1653), .A(N1592), .B(N1588));
AO21XL inst_cellmath__201_0_I874 (.Y(N1654), .A0(N1594), .A1(N1589), .B0(N1593));
AND2XL inst_cellmath__201_0_I875 (.Y(N1655), .A(N1594), .B(N1590));
AO21XL inst_cellmath__201_0_I876 (.Y(N1656), .A0(N1596), .A1(N1591), .B0(N1595));
AND2XL inst_cellmath__201_0_I877 (.Y(N1657), .A(N1596), .B(N1592));
AO21XL inst_cellmath__201_0_I878 (.Y(N1658), .A0(N1598), .A1(N1593), .B0(N1597));
AND2XL inst_cellmath__201_0_I879 (.Y(N1659), .A(N1598), .B(N1594));
AO21XL inst_cellmath__201_0_I880 (.Y(N1660), .A0(N1600), .A1(N1595), .B0(N1599));
AND2XL inst_cellmath__201_0_I881 (.Y(N1661), .A(N1600), .B(N1596));
AO21XL inst_cellmath__201_0_I882 (.Y(N1662), .A0(N1602), .A1(N1597), .B0(N1601));
AND2XL inst_cellmath__201_0_I883 (.Y(N1663), .A(N1602), .B(N1598));
AO21XL inst_cellmath__201_0_I884 (.Y(N1664), .A0(N1604), .A1(N1599), .B0(N1603));
AND2XL inst_cellmath__201_0_I885 (.Y(N1665), .A(N1604), .B(N1600));
AO21XL inst_cellmath__201_0_I886 (.Y(N1666), .A0(N1606), .A1(N1601), .B0(N1605));
AND2XL inst_cellmath__201_0_I887 (.Y(N1667), .A(N1606), .B(N1602));
AO21XL inst_cellmath__201_0_I888 (.Y(N1668), .A0(N1608), .A1(N1603), .B0(N1607));
AND2XL inst_cellmath__201_0_I889 (.Y(N1669), .A(N1608), .B(N1604));
AO21XL inst_cellmath__201_0_I890 (.Y(N1670), .A0(N1610), .A1(N1605), .B0(N1609));
AND2XL inst_cellmath__201_0_I891 (.Y(N1671), .A(N1610), .B(N1606));
AO21XL inst_cellmath__201_0_I892 (.Y(N1672), .A0(N1612), .A1(N1607), .B0(N1611));
AND2XL inst_cellmath__201_0_I893 (.Y(N1673), .A(N1612), .B(N1608));
AO21XL inst_cellmath__201_0_I894 (.Y(N1674), .A0(N1614), .A1(N1609), .B0(N1613));
AND2XL inst_cellmath__201_0_I895 (.Y(N1675), .A(N1614), .B(N1610));
AO21XL inst_cellmath__201_0_I896 (.Y(N1676), .A0(N1616), .A1(N1611), .B0(N1615));
AND2XL inst_cellmath__201_0_I897 (.Y(N1677), .A(N1616), .B(N1612));
AO21XL inst_cellmath__201_0_I898 (.Y(N1678), .A0(N1618), .A1(N1613), .B0(N1617));
AND2XL inst_cellmath__201_0_I899 (.Y(N1679), .A(N1618), .B(N1614));
AO21XL inst_cellmath__201_0_I900 (.Y(N1680), .A0(N1620), .A1(N1615), .B0(N1619));
AND2XL inst_cellmath__201_0_I901 (.Y(N1681), .A(N1620), .B(N1616));
AO21XL inst_cellmath__201_0_I902 (.Y(N1682), .A0(N1622), .A1(N1617), .B0(N1621));
AND2XL inst_cellmath__201_0_I903 (.Y(N1683), .A(N1622), .B(N1618));
AO21XL inst_cellmath__201_0_I904 (.Y(N1684), .A0(N1624), .A1(N1619), .B0(N1623));
AND2XL inst_cellmath__201_0_I905 (.Y(N1685), .A(N1624), .B(N1620));
AO21XL inst_cellmath__201_0_I906 (.Y(N1686), .A0(N1626), .A1(N1621), .B0(N1625));
AND2XL inst_cellmath__201_0_I907 (.Y(N1687), .A(N1626), .B(N1622));
AO21XL inst_cellmath__201_0_I908 (.Y(N1688), .A0(N1628), .A1(N1623), .B0(N1627));
AND2XL inst_cellmath__201_0_I909 (.Y(N1689), .A(N1628), .B(N1624));
AO21XL inst_cellmath__201_0_I910 (.Y(N1690), .A0(N1630), .A1(N1625), .B0(N1629));
AND2XL inst_cellmath__201_0_I911 (.Y(N1691), .A(N1630), .B(N1626));
AO21XL inst_cellmath__201_0_I912 (.Y(N1692), .A0(N1632), .A1(N1627), .B0(N1631));
AND2XL inst_cellmath__201_0_I913 (.Y(N1693), .A(N1632), .B(N1628));
AO21XL inst_cellmath__201_0_I914 (.Y(N1694), .A0(N1634), .A1(N1629), .B0(N1633));
AND2XL inst_cellmath__201_0_I915 (.Y(N1695), .A(N1634), .B(N1630));
AO21XL inst_cellmath__201_0_I916 (.Y(N1696), .A0(N1636), .A1(N1631), .B0(N1635));
AND2XL inst_cellmath__201_0_I917 (.Y(N1697), .A(N1636), .B(N1632));
AO21XL inst_cellmath__201_0_I918 (.Y(N1698), .A0(N1638), .A1(N1633), .B0(N1637));
AND2XL inst_cellmath__201_0_I919 (.Y(N1699), .A(N1638), .B(N1634));
AO21XL inst_cellmath__201_0_I920 (.Y(N1700), .A0(N1640), .A1(N1635), .B0(N1639));
AND2XL inst_cellmath__201_0_I921 (.Y(N1701), .A(N1640), .B(N1636));
AO22XL inst_cellmath__201_0_I1299 (.Y(N1702), .A0(N1049), .A1(N1580), .B0(N1643), .B1(N1637));
AND2XL inst_cellmath__201_0_I923 (.Y(N1703), .A(N1643), .B(N1638));
AO21XL inst_cellmath__201_0_I932 (.Y(N1712), .A0(N1653), .A1(N1524), .B0(N1652));
AO21XL inst_cellmath__201_0_I934 (.Y(N1714), .A0(N1655), .A1(N1585), .B0(N1654));
AO21XL inst_cellmath__201_0_I936 (.Y(N1716), .A0(N1657), .A1(N1648), .B0(N1656));
AO21XL inst_cellmath__201_0_I938 (.Y(N1718), .A0(N1659), .A1(N1650), .B0(N1658));
AO21XL inst_cellmath__201_0_I940 (.Y(N1720), .A0(N1661), .A1(N1652), .B0(N1660));
AND2XL inst_cellmath__201_0_I941 (.Y(N1721), .A(N1661), .B(N1653));
AO21XL inst_cellmath__201_0_I942 (.Y(N1722), .A0(N1663), .A1(N1654), .B0(N1662));
AND2XL inst_cellmath__201_0_I943 (.Y(N1723), .A(N1663), .B(N1655));
AO21XL inst_cellmath__201_0_I944 (.Y(N1724), .A0(N1665), .A1(N1656), .B0(N1664));
AND2XL inst_cellmath__201_0_I945 (.Y(N1725), .A(N1665), .B(N1657));
AO21XL inst_cellmath__201_0_I946 (.Y(N1726), .A0(N1667), .A1(N1658), .B0(N1666));
AND2XL inst_cellmath__201_0_I947 (.Y(N1727), .A(N1667), .B(N1659));
AO21XL inst_cellmath__201_0_I948 (.Y(N1728), .A0(N1669), .A1(N1660), .B0(N1668));
AND2XL inst_cellmath__201_0_I949 (.Y(N1729), .A(N1669), .B(N1661));
AO21XL inst_cellmath__201_0_I950 (.Y(N1730), .A0(N1671), .A1(N1662), .B0(N1670));
AND2XL inst_cellmath__201_0_I951 (.Y(N1731), .A(N1671), .B(N1663));
AO21XL inst_cellmath__201_0_I952 (.Y(N1732), .A0(N1673), .A1(N1664), .B0(N1672));
AND2XL inst_cellmath__201_0_I953 (.Y(N1733), .A(N1673), .B(N1665));
AO21XL inst_cellmath__201_0_I954 (.Y(N1734), .A0(N1675), .A1(N1666), .B0(N1674));
AND2XL inst_cellmath__201_0_I955 (.Y(N1735), .A(N1675), .B(N1667));
AO21XL inst_cellmath__201_0_I956 (.Y(N1736), .A0(N1677), .A1(N1668), .B0(N1676));
AND2XL inst_cellmath__201_0_I957 (.Y(N1737), .A(N1677), .B(N1669));
AO21XL inst_cellmath__201_0_I958 (.Y(N1738), .A0(N1679), .A1(N1670), .B0(N1678));
AND2XL inst_cellmath__201_0_I959 (.Y(N1739), .A(N1679), .B(N1671));
AO21XL inst_cellmath__201_0_I960 (.Y(N1740), .A0(N1681), .A1(N1672), .B0(N1680));
AND2XL inst_cellmath__201_0_I961 (.Y(N1741), .A(N1681), .B(N1673));
AO21XL inst_cellmath__201_0_I962 (.Y(N1742), .A0(N1683), .A1(N1674), .B0(N1682));
AND2XL inst_cellmath__201_0_I963 (.Y(N1743), .A(N1683), .B(N1675));
AO21XL inst_cellmath__201_0_I964 (.Y(N1744), .A0(N1685), .A1(N1676), .B0(N1684));
AND2XL inst_cellmath__201_0_I965 (.Y(N1745), .A(N1685), .B(N1677));
AO21XL inst_cellmath__201_0_I966 (.Y(N1746), .A0(N1687), .A1(N1678), .B0(N1686));
AND2XL inst_cellmath__201_0_I967 (.Y(N1747), .A(N1687), .B(N1679));
AO21XL inst_cellmath__201_0_I968 (.Y(N1748), .A0(N1689), .A1(N1680), .B0(N1688));
AND2XL inst_cellmath__201_0_I969 (.Y(N1749), .A(N1689), .B(N1681));
AO21XL inst_cellmath__201_0_I970 (.Y(N1750), .A0(N1691), .A1(N1682), .B0(N1690));
AND2XL inst_cellmath__201_0_I971 (.Y(N1751), .A(N1691), .B(N1683));
AO21XL inst_cellmath__201_0_I972 (.Y(N1752), .A0(N1693), .A1(N1684), .B0(N1692));
AND2XL inst_cellmath__201_0_I973 (.Y(N1753), .A(N1693), .B(N1685));
AO21XL inst_cellmath__201_0_I974 (.Y(N1754), .A0(N1695), .A1(N1686), .B0(N1694));
AND2XL inst_cellmath__201_0_I975 (.Y(N1755), .A(N1695), .B(N1687));
AO21XL inst_cellmath__201_0_I976 (.Y(N1756), .A0(N1697), .A1(N1688), .B0(N1696));
AND2XL inst_cellmath__201_0_I977 (.Y(N1757), .A(N1697), .B(N1689));
AO21XL inst_cellmath__201_0_I978 (.Y(N1758), .A0(N1699), .A1(N1690), .B0(N1698));
AND2XL inst_cellmath__201_0_I979 (.Y(N1759), .A(N1699), .B(N1691));
AO21XL inst_cellmath__201_0_I980 (.Y(N1760), .A0(N1701), .A1(N1692), .B0(N1700));
AND2XL inst_cellmath__201_0_I981 (.Y(N1761), .A(N1701), .B(N1693));
AO21XL inst_cellmath__201_0_I982 (.Y(N1762), .A0(N1703), .A1(N1694), .B0(N1702));
AND2XL inst_cellmath__201_0_I983 (.Y(N1763), .A(N1703), .B(N1695));
AO21XL inst_cellmath__201_0_I1000 (.Y(N1780), .A0(N1721), .A1(N1524), .B0(N1720));
AO21XL inst_cellmath__201_0_I1002 (.Y(N1782), .A0(N1723), .A1(N1585), .B0(N1722));
AO21XL inst_cellmath__201_0_I1004 (.Y(N1784), .A0(N1725), .A1(N1648), .B0(N1724));
AO21XL inst_cellmath__201_0_I1006 (.Y(N1786), .A0(N1727), .A1(N1650), .B0(N1726));
AO21XL inst_cellmath__201_0_I1008 (.Y(N1788), .A0(N1729), .A1(N1712), .B0(N1728));
AO21XL inst_cellmath__201_0_I1010 (.Y(N1790), .A0(N1731), .A1(N1714), .B0(N1730));
AO21XL inst_cellmath__201_0_I1016 (.Y(N1796), .A0(N1737), .A1(N1720), .B0(N1736));
AND2XL inst_cellmath__201_0_I1017 (.Y(N1797), .A(N1737), .B(N1721));
AO21XL inst_cellmath__201_0_I1018 (.Y(N1798), .A0(N1739), .A1(N1722), .B0(N1738));
AND2XL inst_cellmath__201_0_I1019 (.Y(N1799), .A(N1739), .B(N1723));
AO21XL inst_cellmath__201_0_I1020 (.Y(N1800), .A0(N1741), .A1(N1724), .B0(N1740));
AND2XL inst_cellmath__201_0_I1021 (.Y(N1801), .A(N1741), .B(N1725));
AO21XL inst_cellmath__201_0_I1022 (.Y(N1802), .A0(N1743), .A1(N1726), .B0(N1742));
AND2XL inst_cellmath__201_0_I1023 (.Y(N1803), .A(N1743), .B(N1727));
AO21XL inst_cellmath__201_0_I1024 (.Y(N1804), .A0(N1745), .A1(N1728), .B0(N1744));
AND2XL inst_cellmath__201_0_I1025 (.Y(N1805), .A(N1745), .B(N1729));
AO21XL inst_cellmath__201_0_I1026 (.Y(N1806), .A0(N1747), .A1(N1730), .B0(N1746));
AND2XL inst_cellmath__201_0_I1027 (.Y(N1807), .A(N1747), .B(N1731));
AO21XL inst_cellmath__201_0_I1028 (.Y(N1808), .A0(N1749), .A1(N1732), .B0(N1748));
AND2XL inst_cellmath__201_0_I1029 (.Y(N1809), .A(N1749), .B(N1733));
AO21XL inst_cellmath__201_0_I1030 (.Y(N1810), .A0(N1751), .A1(N1734), .B0(N1750));
AND2XL inst_cellmath__201_0_I1031 (.Y(N1811), .A(N1751), .B(N1735));
AO21XL inst_cellmath__201_0_I1032 (.Y(N1812), .A0(N1753), .A1(N1736), .B0(N1752));
AND2XL inst_cellmath__201_0_I1033 (.Y(N1813), .A(N1753), .B(N1737));
AO21XL inst_cellmath__201_0_I1034 (.Y(N1814), .A0(N1755), .A1(N1738), .B0(N1754));
AND2XL inst_cellmath__201_0_I1035 (.Y(N1815), .A(N1755), .B(N1739));
AO21XL inst_cellmath__201_0_I1036 (.Y(N1816), .A0(N1757), .A1(N1740), .B0(N1756));
AND2XL inst_cellmath__201_0_I1037 (.Y(N1817), .A(N1757), .B(N1741));
AO21XL inst_cellmath__201_0_I1038 (.Y(N1818), .A0(N1759), .A1(N1742), .B0(N1758));
AND2XL inst_cellmath__201_0_I1039 (.Y(N1819), .A(N1759), .B(N1743));
AO21XL inst_cellmath__201_0_I1040 (.Y(N1820), .A0(N1761), .A1(N1744), .B0(N1760));
AND2XL inst_cellmath__201_0_I1041 (.Y(N1821), .A(N1761), .B(N1745));
AO21XL inst_cellmath__201_0_I1042 (.Y(N1822), .A0(N1763), .A1(N1746), .B0(N1762));
AND2XL inst_cellmath__201_0_I1043 (.Y(N1823), .A(N1763), .B(N1747));
AOI21XL inst_cellmath__201_0_I1591 (.Y(N2440), .A0(N1733), .A1(N1716), .B0(N1732));
AOI21XL inst_cellmath__201_0_I1592 (.Y(N2441), .A0(N1735), .A1(N1718), .B0(N1734));
AO21XL inst_cellmath__201_0_I1076 (.Y(N1856), .A0(N1797), .A1(N1524), .B0(N1796));
AO21XL inst_cellmath__201_0_I1078 (.Y(N1858), .A0(N1799), .A1(N1585), .B0(N1798));
AO21XL inst_cellmath__201_0_I1080 (.Y(N1860), .A0(N1801), .A1(N1648), .B0(N1800));
AO21XL inst_cellmath__201_0_I1082 (.Y(N1862), .A0(N1803), .A1(N1650), .B0(N1802));
AO21XL inst_cellmath__201_0_I1084 (.Y(N1864), .A0(N1805), .A1(N1712), .B0(N1804));
AO21XL inst_cellmath__201_0_I1086 (.Y(N1866), .A0(N1807), .A1(N1714), .B0(N1806));
AO21XL inst_cellmath__201_0_I1088 (.Y(N1868), .A0(N1809), .A1(N1716), .B0(N1808));
AO21XL inst_cellmath__201_0_I1090 (.Y(N1870), .A0(N1811), .A1(N1718), .B0(N1810));
AO21XL inst_cellmath__201_0_I1092 (.Y(N1872), .A0(N1813), .A1(N1780), .B0(N1812));
AO21XL inst_cellmath__201_0_I1094 (.Y(N1874), .A0(N1815), .A1(N1782), .B0(N1814));
AO21XL inst_cellmath__201_0_I1096 (.Y(N1876), .A0(N1817), .A1(N1784), .B0(N1816));
AO21XL inst_cellmath__201_0_I1098 (.Y(N1878), .A0(N1819), .A1(N1786), .B0(N1818));
AO21XL inst_cellmath__201_0_I1100 (.Y(N1880), .A0(N1821), .A1(N1788), .B0(N1820));
AO21XL inst_cellmath__201_0_I1102 (.Y(inst_cellmath__201_0_out0[49]), .A0(N1823), .A1(N1790), .B0(N1822));
NAND2BXL inst_cellmath__201_0_I1109 (.Y(N1889), .AN(N1526), .B(N1527));
NAND2BXL inst_cellmath__201_0_I1112 (.Y(N1892), .AN(N1528), .B(N1529));
NAND2BXL inst_cellmath__201_0_I1115 (.Y(N1895), .AN(N1530), .B(N1531));
NAND2BXL inst_cellmath__201_0_I1118 (.Y(N1898), .AN(N1532), .B(N1533));
NAND2BXL inst_cellmath__201_0_I1121 (.Y(N1901), .AN(N1534), .B(N1535));
NAND2BXL inst_cellmath__201_0_I1124 (.Y(N1904), .AN(N1536), .B(N1537));
NAND2BXL inst_cellmath__201_0_I1127 (.Y(N1907), .AN(N1538), .B(N1539));
NAND2BXL inst_cellmath__201_0_I1130 (.Y(N1910), .AN(N1540), .B(N1541));
NAND2BXL inst_cellmath__201_0_I1133 (.Y(N1913), .AN(N1542), .B(N1543));
NAND2BXL inst_cellmath__201_0_I1136 (.Y(N1916), .AN(N1544), .B(N1545));
NAND2BXL inst_cellmath__201_0_I1139 (.Y(N1919), .AN(N1546), .B(N1547));
NAND2BXL inst_cellmath__201_0_I1142 (.Y(N1922), .AN(N1548), .B(N1549));
NAND2BXL inst_cellmath__201_0_I1145 (.Y(N1925), .AN(N1550), .B(N1551));
NAND2BXL inst_cellmath__201_0_I1148 (.Y(N1928), .AN(N1552), .B(N1553));
NAND2BXL inst_cellmath__201_0_I1151 (.Y(N1931), .AN(N1554), .B(N1555));
NAND2BXL inst_cellmath__201_0_I1154 (.Y(N1934), .AN(N1556), .B(N1557));
NAND2BXL inst_cellmath__201_0_I1157 (.Y(N1937), .AN(N1558), .B(N1559));
NAND2BXL inst_cellmath__201_0_I1160 (.Y(N1940), .AN(N1560), .B(N1561));
NAND2BXL inst_cellmath__201_0_I1163 (.Y(N1943), .AN(N1562), .B(N1563));
NAND2BXL inst_cellmath__201_0_I1166 (.Y(N1946), .AN(N1564), .B(N1565));
NAND2BXL inst_cellmath__201_0_I1169 (.Y(N1949), .AN(N1566), .B(N1567));
NAND2BXL inst_cellmath__201_0_I1172 (.Y(N1952), .AN(N1568), .B(N1569));
NAND2BXL inst_cellmath__201_0_I1175 (.Y(N1955), .AN(N1570), .B(N1571));
NAND2BXL inst_cellmath__201_0_I1178 (.Y(N1958), .AN(N1572), .B(N1573));
NAND2BXL inst_cellmath__201_0_I1181 (.Y(N1961), .AN(N1574), .B(N1575));
NAND2BXL inst_cellmath__201_0_I1184 (.Y(N1964), .AN(N1576), .B(N1577));
NAND2BXL inst_cellmath__201_0_I1187 (.Y(N1967), .AN(N1578), .B(N1579));
NAND2BXL inst_cellmath__201_0_I1190 (.Y(N1970), .AN(N1580), .B(N1581));
XOR2XL inst_cellmath__201_0_I1593 (.Y(inst_cellmath__201_0_out0[20]), .A(N1524), .B(N1889));
XOR2XL inst_cellmath__201_0_I1594 (.Y(inst_cellmath__201_0_out0[21]), .A(N1585), .B(N1892));
XOR2XL inst_cellmath__201_0_I1595 (.Y(inst_cellmath__201_0_out0[22]), .A(N1648), .B(N1895));
XOR2XL inst_cellmath__201_0_I1596 (.Y(inst_cellmath__201_0_out0[23]), .A(N1650), .B(N1898));
XOR2XL inst_cellmath__201_0_I1597 (.Y(inst_cellmath__201_0_out0[24]), .A(N1712), .B(N1901));
XOR2XL inst_cellmath__201_0_I1598 (.Y(inst_cellmath__201_0_out0[25]), .A(N1714), .B(N1904));
XOR2XL inst_cellmath__201_0_I1599 (.Y(inst_cellmath__201_0_out0[26]), .A(N1716), .B(N1907));
XOR2XL inst_cellmath__201_0_I1600 (.Y(inst_cellmath__201_0_out0[27]), .A(N1718), .B(N1910));
XOR2XL inst_cellmath__201_0_I1601 (.Y(inst_cellmath__201_0_out0[28]), .A(N1780), .B(N1913));
XOR2XL inst_cellmath__201_0_I1602 (.Y(inst_cellmath__201_0_out0[29]), .A(N1782), .B(N1916));
XOR2XL inst_cellmath__201_0_I1603 (.Y(inst_cellmath__201_0_out0[30]), .A(N1784), .B(N1919));
XOR2XL inst_cellmath__201_0_I1604 (.Y(inst_cellmath__201_0_out0[31]), .A(N1786), .B(N1922));
XOR2XL inst_cellmath__201_0_I1605 (.Y(inst_cellmath__201_0_out0[32]), .A(N1788), .B(N1925));
XOR2XL inst_cellmath__201_0_I1606 (.Y(inst_cellmath__201_0_out0[33]), .A(N1790), .B(N1928));
XNOR2X1 inst_cellmath__201_0_I1209 (.Y(inst_cellmath__201_0_out0[34]), .A(N2440), .B(N1931));
XNOR2X1 inst_cellmath__201_0_I1210 (.Y(inst_cellmath__201_0_out0[35]), .A(N2441), .B(N1934));
XOR2XL inst_cellmath__201_0_I1211 (.Y(inst_cellmath__201_0_out0[36]), .A(N1856), .B(N1937));
XOR2XL inst_cellmath__201_0_I1212 (.Y(inst_cellmath__201_0_out0[37]), .A(N1858), .B(N1940));
XOR2XL inst_cellmath__201_0_I1213 (.Y(inst_cellmath__201_0_out0[38]), .A(N1860), .B(N1943));
XOR2XL inst_cellmath__201_0_I1214 (.Y(inst_cellmath__201_0_out0[39]), .A(N1862), .B(N1946));
XOR2XL inst_cellmath__201_0_I1215 (.Y(inst_cellmath__201_0_out0[40]), .A(N1864), .B(N1949));
XOR2XL inst_cellmath__201_0_I1216 (.Y(inst_cellmath__201_0_out0[41]), .A(N1866), .B(N1952));
XOR2XL inst_cellmath__201_0_I1217 (.Y(inst_cellmath__201_0_out0[42]), .A(N1868), .B(N1955));
XOR2XL inst_cellmath__201_0_I1218 (.Y(inst_cellmath__201_0_out0[43]), .A(N1870), .B(N1958));
XOR2XL inst_cellmath__201_0_I1219 (.Y(inst_cellmath__201_0_out0[44]), .A(N1872), .B(N1961));
XOR2XL inst_cellmath__201_0_I1220 (.Y(inst_cellmath__201_0_out0[45]), .A(N1874), .B(N1964));
XOR2XL inst_cellmath__201_0_I1221 (.Y(inst_cellmath__201_0_out0[46]), .A(N1876), .B(N1967));
XOR2XL inst_cellmath__201_0_I1222 (.Y(inst_cellmath__201_0_out0[47]), .A(N1878), .B(N1970));
XNOR2X1 inst_cellmath__201_0_I1223 (.Y(inst_cellmath__201_0_out0[48]), .A(N1880), .B(N1049));
assign inst_cellmath__203__W1[0] = inst_cellmath__201_0_in1[0];
assign inst_cellmath__203__W1[1] = inst_cellmath__201_0_in0[1];
assign inst_cellmath__203__W1[2] = inst_cellmath__201_0_in0[2];
assign inst_cellmath__203__W1[3] = inst_cellmath__201_0_in0[3];
assign inst_cellmath__203__W1[4] = inst_cellmath__201_0_in0[4];
assign inst_cellmath__203__W1[5] = inst_cellmath__201_0_in0[5];
assign inst_cellmath__203__W1[6] = inst_cellmath__201_0_in0[6];
assign inst_cellmath__203__W1[7] = inst_cellmath__201_0_in0[7];
assign inst_cellmath__203__W1[8] = inst_cellmath__201_0_in0[8];
assign inst_cellmath__203__W1[9] = inst_cellmath__201_0_in0[9];
assign inst_cellmath__203__W1[10] = inst_cellmath__201_0_in0[10];
assign inst_cellmath__203__W1[11] = inst_cellmath__201_0_in0[11];
assign inst_cellmath__203__W1[12] = inst_cellmath__201_0_in0[12];
assign inst_cellmath__203__W1[13] = inst_cellmath__201_0_in0[13];
assign inst_cellmath__203__W1[14] = inst_cellmath__201_0_in0[14];
assign inst_cellmath__203__W1[15] = inst_cellmath__201_0_in0[15];
assign inst_cellmath__203__W1[16] = inst_cellmath__201_0_in0[16];
assign inst_cellmath__203__W1[17] = inst_cellmath__201_0_in0[17];
assign inst_cellmath__203__W1[18] = inst_cellmath__201_0_in0[18];
assign inst_cellmath__203__W1[19] = inst_cellmath__201_0_in0[19];
assign inst_cellmath__203__W1[20] = inst_cellmath__201_0_in0[20];
assign inst_cellmath__203__W1[21] = inst_cellmath__201_0_in0[21];
assign inst_cellmath__203__W1[22] = inst_cellmath__201_0_in0[22];
assign inst_cellmath__203__W1[23] = inst_cellmath__201_0_in0[23];
assign inst_cellmath__203__W1[24] = inst_cellmath__201_0_in0[24];
assign inst_cellmath__203__W1[25] = inst_cellmath__201_0_in0[25];
assign inst_cellmath__203__W1[26] = inst_cellmath__201_0_in0[26];
assign inst_cellmath__203__W1[27] = inst_cellmath__201_0_in0[27];
assign inst_cellmath__203__W1[28] = inst_cellmath__201_0_in0[28];
assign inst_cellmath__203__W1[29] = inst_cellmath__201_0_in0[29];
assign inst_cellmath__203__W1[30] = inst_cellmath__201_0_in0[30];
assign inst_cellmath__203__W1[31] = inst_cellmath__201_0_in0[31];
assign inst_cellmath__203__W1[32] = inst_cellmath__201_0_in0[32];
assign inst_cellmath__203__W1[33] = inst_cellmath__201_0_in1[33];
assign inst_cellmath__203__W1[34] = inst_cellmath__201_0_in0[34];
assign inst_cellmath__203__W1[35] = inst_cellmath__201_0_in1[35];
assign inst_cellmath__203__W1[36] = inst_cellmath__201_0_in0[36];
assign inst_cellmath__203__W1[37] = inst_cellmath__201_0_in0[37];
assign inst_cellmath__203__W1[38] = inst_cellmath__201_0_in0[38];
assign inst_cellmath__203__W1[39] = inst_cellmath__201_0_in0[39];
assign inst_cellmath__203__W1[40] = inst_cellmath__201_0_in0[40];
assign inst_cellmath__203__W1[41] = inst_cellmath__201_0_in0[41];
assign inst_cellmath__203__W1[42] = inst_cellmath__201_0_in0[42];
assign inst_cellmath__203__W1[43] = inst_cellmath__201_0_in0[43];
assign inst_cellmath__203__W1[44] = inst_cellmath__201_0_in0[44];
assign inst_cellmath__203__W1[45] = inst_cellmath__201_0_in0[45];
endmodule

module cynw_cm_float_cos_inst_cellmath__200_0_bdw1114505291_bdw (
	inst_cellmath__200_0_out0,
	inst_cellmath__200_0_in0
	); /* architecture "gate_level" */ 
output [48:0] inst_cellmath__200_0_out0;
input [49:0] inst_cellmath__200_0_in0;
wire N202;
BUFX2 inst_cellmath__200_0_I52 (.Y(N202), .A(inst_cellmath__200_0_in0[49]));
NOR2BX1 inst_cellmath__200_0_I0 (.Y(inst_cellmath__200_0_out0[0]), .AN(inst_cellmath__200_0_in0[0]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I1 (.Y(inst_cellmath__200_0_out0[1]), .AN(inst_cellmath__200_0_in0[1]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I2 (.Y(inst_cellmath__200_0_out0[2]), .AN(inst_cellmath__200_0_in0[2]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I3 (.Y(inst_cellmath__200_0_out0[3]), .AN(inst_cellmath__200_0_in0[3]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I4 (.Y(inst_cellmath__200_0_out0[4]), .AN(inst_cellmath__200_0_in0[4]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I5 (.Y(inst_cellmath__200_0_out0[5]), .AN(inst_cellmath__200_0_in0[5]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I6 (.Y(inst_cellmath__200_0_out0[6]), .AN(inst_cellmath__200_0_in0[6]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I7 (.Y(inst_cellmath__200_0_out0[7]), .AN(inst_cellmath__200_0_in0[7]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I8 (.Y(inst_cellmath__200_0_out0[8]), .AN(inst_cellmath__200_0_in0[8]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I9 (.Y(inst_cellmath__200_0_out0[9]), .AN(inst_cellmath__200_0_in0[9]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I10 (.Y(inst_cellmath__200_0_out0[10]), .AN(inst_cellmath__200_0_in0[10]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I11 (.Y(inst_cellmath__200_0_out0[11]), .AN(inst_cellmath__200_0_in0[11]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I12 (.Y(inst_cellmath__200_0_out0[12]), .AN(inst_cellmath__200_0_in0[12]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I13 (.Y(inst_cellmath__200_0_out0[13]), .AN(inst_cellmath__200_0_in0[13]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I14 (.Y(inst_cellmath__200_0_out0[14]), .AN(inst_cellmath__200_0_in0[14]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I15 (.Y(inst_cellmath__200_0_out0[15]), .AN(inst_cellmath__200_0_in0[15]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I16 (.Y(inst_cellmath__200_0_out0[16]), .AN(inst_cellmath__200_0_in0[16]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I17 (.Y(inst_cellmath__200_0_out0[17]), .AN(inst_cellmath__200_0_in0[17]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I18 (.Y(inst_cellmath__200_0_out0[18]), .AN(inst_cellmath__200_0_in0[18]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I19 (.Y(inst_cellmath__200_0_out0[19]), .AN(inst_cellmath__200_0_in0[19]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I20 (.Y(inst_cellmath__200_0_out0[20]), .AN(inst_cellmath__200_0_in0[20]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I21 (.Y(inst_cellmath__200_0_out0[21]), .AN(inst_cellmath__200_0_in0[21]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I22 (.Y(inst_cellmath__200_0_out0[22]), .AN(inst_cellmath__200_0_in0[22]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I23 (.Y(inst_cellmath__200_0_out0[23]), .AN(inst_cellmath__200_0_in0[23]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I24 (.Y(inst_cellmath__200_0_out0[24]), .AN(inst_cellmath__200_0_in0[24]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I25 (.Y(inst_cellmath__200_0_out0[25]), .AN(inst_cellmath__200_0_in0[25]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I26 (.Y(inst_cellmath__200_0_out0[26]), .AN(inst_cellmath__200_0_in0[26]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I27 (.Y(inst_cellmath__200_0_out0[27]), .AN(inst_cellmath__200_0_in0[27]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I28 (.Y(inst_cellmath__200_0_out0[28]), .AN(inst_cellmath__200_0_in0[28]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I29 (.Y(inst_cellmath__200_0_out0[29]), .AN(inst_cellmath__200_0_in0[29]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I30 (.Y(inst_cellmath__200_0_out0[30]), .AN(inst_cellmath__200_0_in0[30]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I31 (.Y(inst_cellmath__200_0_out0[31]), .AN(inst_cellmath__200_0_in0[31]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I32 (.Y(inst_cellmath__200_0_out0[32]), .AN(inst_cellmath__200_0_in0[32]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I33 (.Y(inst_cellmath__200_0_out0[33]), .AN(inst_cellmath__200_0_in0[33]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I34 (.Y(inst_cellmath__200_0_out0[34]), .AN(inst_cellmath__200_0_in0[34]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I35 (.Y(inst_cellmath__200_0_out0[35]), .AN(inst_cellmath__200_0_in0[35]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I36 (.Y(inst_cellmath__200_0_out0[36]), .AN(inst_cellmath__200_0_in0[36]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I37 (.Y(inst_cellmath__200_0_out0[37]), .AN(inst_cellmath__200_0_in0[37]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I38 (.Y(inst_cellmath__200_0_out0[38]), .AN(inst_cellmath__200_0_in0[38]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I39 (.Y(inst_cellmath__200_0_out0[39]), .AN(inst_cellmath__200_0_in0[39]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I40 (.Y(inst_cellmath__200_0_out0[40]), .AN(inst_cellmath__200_0_in0[40]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I41 (.Y(inst_cellmath__200_0_out0[41]), .AN(inst_cellmath__200_0_in0[41]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I42 (.Y(inst_cellmath__200_0_out0[42]), .AN(inst_cellmath__200_0_in0[42]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I43 (.Y(inst_cellmath__200_0_out0[43]), .AN(inst_cellmath__200_0_in0[43]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I44 (.Y(inst_cellmath__200_0_out0[44]), .AN(inst_cellmath__200_0_in0[44]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I45 (.Y(inst_cellmath__200_0_out0[45]), .AN(inst_cellmath__200_0_in0[45]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I46 (.Y(inst_cellmath__200_0_out0[46]), .AN(inst_cellmath__200_0_in0[46]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I47 (.Y(inst_cellmath__200_0_out0[47]), .AN(inst_cellmath__200_0_in0[47]), .B(N202));
NOR2BX1 inst_cellmath__200_0_I48 (.Y(inst_cellmath__200_0_out0[48]), .AN(inst_cellmath__200_0_in0[48]), .B(N202));
endmodule

module cynw_cm_float_cos_inst_cellmath__17_0_bdw1114505291_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[0]));
NOR2XL inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[6]), .B(inst_cellmath__17_0_in0[5]));
NOR2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[4]), .B(inst_cellmath__17_0_in0[3]));
NOR2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[2]), .B(inst_cellmath__17_0_in0[1]));
NAND2XL inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_cos_inst_cellmath__46__15__bdw1114505291_bdw (
	inst_cellmath__46__15__out0,
	inst_cellmath__46__15__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__46__15__out0;
input [7:6] inst_cellmath__46__15__in0;
OR2XL inst_cellmath__46__15__I0 (.Y(inst_cellmath__46__15__out0[0]), .A(inst_cellmath__46__15__in0[7]), .B(inst_cellmath__46__15__in0[6]));
endmodule

module cynw_cm_float_cos_inst_cellmath__46_0_bdw1114505291_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__46_0_out0;
input [0:0] inst_cellmath__46_0_in0;
input [8:8] inst_cellmath__46_0_in1;
NOR2BX1 inst_cellmath__46_0_I3 (.Y(inst_cellmath__46_0_out0), .AN(inst_cellmath__46_0_in0[0]), .B(inst_cellmath__46_0_in1[8]));
endmodule

module cynw_cm_float_cos_inst_cellmath__21_0_bdw1114505291_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input [7:0] inst_cellmath__21_0_in0;
wire N66,N70;
AOI211XL inst_cellmath__21_0_I39 (.Y(N66), .A0(inst_cellmath__21_0_in0[2]), .A1(inst_cellmath__21_0_in0[1]), .B0(inst_cellmath__21_0_in0[3]), .C0(inst_cellmath__21_0_in0[4]));
NAND3BXL inst_cellmath__21_0_I37 (.Y(N70), .AN(N66), .B(inst_cellmath__21_0_in0[5]), .C(inst_cellmath__21_0_in0[6]));
NOR2BX1 inst_cellmath__21_0_I38 (.Y(inst_cellmath__21_0_out0), .AN(N70), .B(inst_cellmath__21_0_in0[7]));
endmodule

module cynw_cm_float_cos_inst_cellmath__83__62__bdw1114505291_bdw (
	inst_cellmath__83__62__out0,
	inst_cellmath__83__62__in0,
	inst_cellmath__83__62__in1,
	inst_cellmath__83__62__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__83__62__out0;
input  inst_cellmath__83__62__in0,
	inst_cellmath__83__62__in1,
	inst_cellmath__83__62__in2;
OR3XL inst_cellmath__83__62__I4 (.Y(inst_cellmath__83__62__out0[0]), .A(inst_cellmath__83__62__in2), .B(inst_cellmath__83__62__in1), .C(inst_cellmath__83__62__in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__19_0_bdw1114505291_bdw (
	inst_cellmath__19_0_out0,
	inst_cellmath__19_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19_0_out0;
input [7:0] inst_cellmath__19_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__19_0_I0 (.Y(N11), .A(inst_cellmath__19_0_in0[7]), .B(inst_cellmath__19_0_in0[0]));
NAND2XL inst_cellmath__19_0_I1 (.Y(N12), .A(inst_cellmath__19_0_in0[6]), .B(inst_cellmath__19_0_in0[5]));
NAND2XL inst_cellmath__19_0_I2 (.Y(N13), .A(inst_cellmath__19_0_in0[4]), .B(inst_cellmath__19_0_in0[3]));
NAND2XL inst_cellmath__19_0_I3 (.Y(N14), .A(inst_cellmath__19_0_in0[2]), .B(inst_cellmath__19_0_in0[1]));
NOR2XL inst_cellmath__19_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__19_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__19_0_I6 (.Y(inst_cellmath__19_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_cos_inst_cellmath__24_0_bdw1114505291_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__24_0_I1 (.Y(N27), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
NOR2XL inst_cellmath__24_0_I2 (.Y(N28), .A(inst_cellmath__24_0_in0[20]), .B(inst_cellmath__24_0_in0[19]));
NOR2XL inst_cellmath__24_0_I3 (.Y(N29), .A(inst_cellmath__24_0_in0[18]), .B(inst_cellmath__24_0_in0[17]));
NOR2XL inst_cellmath__24_0_I4 (.Y(N30), .A(inst_cellmath__24_0_in0[16]), .B(inst_cellmath__24_0_in0[15]));
NOR2XL inst_cellmath__24_0_I5 (.Y(N31), .A(inst_cellmath__24_0_in0[14]), .B(inst_cellmath__24_0_in0[13]));
NOR2XL inst_cellmath__24_0_I6 (.Y(N32), .A(inst_cellmath__24_0_in0[12]), .B(inst_cellmath__24_0_in0[11]));
NOR2XL inst_cellmath__24_0_I7 (.Y(N33), .A(inst_cellmath__24_0_in0[10]), .B(inst_cellmath__24_0_in0[9]));
NOR2XL inst_cellmath__24_0_I8 (.Y(N34), .A(inst_cellmath__24_0_in0[8]), .B(inst_cellmath__24_0_in0[7]));
NOR2XL inst_cellmath__24_0_I9 (.Y(N35), .A(inst_cellmath__24_0_in0[6]), .B(inst_cellmath__24_0_in0[5]));
NOR2XL inst_cellmath__24_0_I10 (.Y(N36), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in0[3]));
NAND2XL inst_cellmath__24_0_I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__24_0_I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__24_0_I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__24_0_I25 (.Y(N44), .A(inst_cellmath__24_0_in0[0]), .B(inst_cellmath__24_0_in0[1]), .C(inst_cellmath__24_0_in0[2]), .D(N39));
NOR2XL inst_cellmath__24_0_I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__24_0_I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__24_0_I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__24_0_I23 (.Y(inst_cellmath__24_0_out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_cos_inst_cellmath__69_0_bdw1114505291_bdw (
	inst_cellmath__69_0_out0,
	inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__69_0_out0;
input  inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1;
NOR2BX1 inst_cellmath__69_0_I2 (.Y(inst_cellmath__69_0_out0), .AN(inst_cellmath__69_0_in1), .B(inst_cellmath__69_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__82_0_bdw1114505291_bdw (
	inst_cellmath__82_0_out0,
	inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__82_0_out0;
input  inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1;
OR2XL inst_cellmath__82_0_I0 (.Y(inst_cellmath__82_0_out0), .A(inst_cellmath__82_0_in1), .B(inst_cellmath__82_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__66_0_bdw1114505291_bdw (
	inst_cellmath__66_0_out0,
	inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__66_0_out0;
input  inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2;
wire N18;
NAND2XL inst_cellmath__66_0_I7 (.Y(N18), .A(inst_cellmath__66_0_in1), .B(inst_cellmath__66_0_in0));
NOR2XL inst_cellmath__66_0_I8 (.Y(inst_cellmath__66_0_out0), .A(inst_cellmath__66_0_in2), .B(N18));
endmodule

module cynw_cm_float_cos_inst_cellmath__67_0_bdw1114505291_bdw (
	inst_cellmath__67_0_out0,
	inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__67_0_out0;
input  inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2;
AND3XL inst_cellmath__67_0_I4 (.Y(inst_cellmath__67_0_out0), .A(inst_cellmath__67_0_in2), .B(inst_cellmath__67_0_in1), .C(inst_cellmath__67_0_in0));
endmodule

module cynw_cm_float_cos_inst_cellmath__68_0_bdw1114505291_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__68_0_out0;
input  inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1;
OR2XL inst_cellmath__68_0_I0 (.Y(inst_cellmath__68_0_out0), .A(inst_cellmath__68_0_in0), .B(inst_cellmath__68_0_in1));
endmodule

module cynw_cm_float_cos_inst_cellmath__228__231__bdw1114505291_bdw (
	inst_cellmath__228__231__out0,
	inst_cellmath__228__231__in0,
	inst_cellmath__228__231__in1,
	inst_cellmath__228__231__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__228__231__out0;
input [0:0] inst_cellmath__228__231__in0;
input  inst_cellmath__228__231__in1,
	inst_cellmath__228__231__in2;
OR3XL inst_cellmath__228__231__I4 (.Y(inst_cellmath__228__231__out0[0]), .A(inst_cellmath__228__231__in1), .B(inst_cellmath__228__231__in2), .C(inst_cellmath__228__231__in0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__219_0_bdw1114505291_bdw (
	inst_cellmath__219_0_out0,
	inst_cellmath__219_0_in0,
	inst_cellmath__219_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__219_0_out0;
input [22:22] inst_cellmath__219_0_in0;
input [48:48] inst_cellmath__219_0_in1;
AND2XL inst_cellmath__219_0_I0 (.Y(inst_cellmath__219_0_out0), .A(inst_cellmath__219_0_in0[22]), .B(inst_cellmath__219_0_in1[48]));
endmodule

module cynw_cm_float_cos_inst_cellmath__211__182__bdw1114505291_bdw (
	inst_cellmath__211__182__out0,
	inst_cellmath__211__182__in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__211__182__out0;
input [47:25] inst_cellmath__211__182__in0;
wire N100,N106,N108,N109,N113,N114,N115 
	,N116,N117,N119,N120,N121,N122,N123,N125 
	,N126,N127,N128,N129,N131,N132,N133,N134 
	,N135,N137,N139,N140,N141,N155,N157,N158 
	,N160,N162,N163,N164,N165,N166,N168,N171 
	,N172,N180,N182,N183,N189,N191,N194,N216 
	,N218,N232,N234,N240,N242;
INVXL inst_cellmath__211__182__I7 (.Y(N100), .A(inst_cellmath__211__182__in0[47]));
INVXL inst_cellmath__211__182__I11 (.Y(N106), .A(inst_cellmath__211__182__in0[25]));
INVXL inst_cellmath__211__182__I12 (.Y(N108), .A(inst_cellmath__211__182__in0[27]));
OAI21XL inst_cellmath__211__182__I13 (.Y(N109), .A0(inst_cellmath__211__182__in0[26]), .A1(N106), .B0(N108));
OR2XL inst_cellmath__211__182__I15 (.Y(N155), .A(inst_cellmath__211__182__in0[27]), .B(inst_cellmath__211__182__in0[26]));
NOR2BX1 inst_cellmath__211__182__I142 (.Y(N113), .AN(inst_cellmath__211__182__in0[28]), .B(inst_cellmath__211__182__in0[29]));
INVXL inst_cellmath__211__182__I18 (.Y(N114), .A(inst_cellmath__211__182__in0[31]));
OAI21XL inst_cellmath__211__182__I19 (.Y(N115), .A0(inst_cellmath__211__182__in0[30]), .A1(N113), .B0(N114));
NOR2XL inst_cellmath__211__182__I20 (.Y(N116), .A(inst_cellmath__211__182__in0[29]), .B(inst_cellmath__211__182__in0[28]));
NOR2XL inst_cellmath__211__182__I21 (.Y(N117), .A(inst_cellmath__211__182__in0[31]), .B(inst_cellmath__211__182__in0[30]));
NOR2BX1 inst_cellmath__211__182__I143 (.Y(N119), .AN(inst_cellmath__211__182__in0[32]), .B(inst_cellmath__211__182__in0[33]));
INVXL inst_cellmath__211__182__I24 (.Y(N120), .A(inst_cellmath__211__182__in0[35]));
OAI21XL inst_cellmath__211__182__I25 (.Y(N121), .A0(inst_cellmath__211__182__in0[34]), .A1(N119), .B0(N120));
NOR2XL inst_cellmath__211__182__I26 (.Y(N122), .A(inst_cellmath__211__182__in0[33]), .B(inst_cellmath__211__182__in0[32]));
NOR2XL inst_cellmath__211__182__I27 (.Y(N123), .A(inst_cellmath__211__182__in0[35]), .B(inst_cellmath__211__182__in0[34]));
NOR2BX1 inst_cellmath__211__182__I144 (.Y(N125), .AN(inst_cellmath__211__182__in0[36]), .B(inst_cellmath__211__182__in0[37]));
INVXL inst_cellmath__211__182__I30 (.Y(N126), .A(inst_cellmath__211__182__in0[39]));
OAI21XL inst_cellmath__211__182__I31 (.Y(N127), .A0(inst_cellmath__211__182__in0[38]), .A1(N125), .B0(N126));
NOR2XL inst_cellmath__211__182__I32 (.Y(N128), .A(inst_cellmath__211__182__in0[37]), .B(inst_cellmath__211__182__in0[36]));
NOR2XL inst_cellmath__211__182__I33 (.Y(N129), .A(inst_cellmath__211__182__in0[39]), .B(inst_cellmath__211__182__in0[38]));
NOR2BX1 inst_cellmath__211__182__I145 (.Y(N131), .AN(inst_cellmath__211__182__in0[40]), .B(inst_cellmath__211__182__in0[41]));
INVXL inst_cellmath__211__182__I36 (.Y(N132), .A(inst_cellmath__211__182__in0[43]));
OAI21XL inst_cellmath__211__182__I37 (.Y(N133), .A0(inst_cellmath__211__182__in0[42]), .A1(N131), .B0(N132));
NOR2XL inst_cellmath__211__182__I38 (.Y(N134), .A(inst_cellmath__211__182__in0[41]), .B(inst_cellmath__211__182__in0[40]));
NOR2XL inst_cellmath__211__182__I39 (.Y(N135), .A(inst_cellmath__211__182__in0[43]), .B(inst_cellmath__211__182__in0[42]));
NOR2BX1 inst_cellmath__211__182__I146 (.Y(N137), .AN(inst_cellmath__211__182__in0[44]), .B(inst_cellmath__211__182__in0[45]));
OAI21XL inst_cellmath__211__182__I43 (.Y(N139), .A0(inst_cellmath__211__182__in0[46]), .A1(N137), .B0(N100));
NOR2XL inst_cellmath__211__182__I44 (.Y(N140), .A(inst_cellmath__211__182__in0[45]), .B(inst_cellmath__211__182__in0[44]));
NOR2XL inst_cellmath__211__182__I45 (.Y(N141), .A(inst_cellmath__211__182__in0[47]), .B(inst_cellmath__211__182__in0[46]));
INVXL inst_cellmath__211__182__I60 (.Y(N157), .A(N117));
AOI21XL inst_cellmath__211__182__I61 (.Y(N158), .A0(N116), .A1(N155), .B0(N157));
NAND2XL inst_cellmath__211__182__I63 (.Y(N160), .A(N117), .B(N116));
NAND2BXL inst_cellmath__211__182__I147 (.Y(N162), .AN(N122), .B(N123));
INVXL inst_cellmath__211__182__I66 (.Y(N163), .A(N129));
AOI21XL inst_cellmath__211__182__I67 (.Y(N164), .A0(N128), .A1(N162), .B0(N163));
NAND2XL inst_cellmath__211__182__I68 (.Y(N165), .A(N123), .B(N122));
NAND2XL inst_cellmath__211__182__I69 (.Y(N166), .A(N129), .B(N128));
NAND2BXL inst_cellmath__211__182__I148 (.Y(N168), .AN(N134), .B(N135));
NAND2XL inst_cellmath__211__182__I74 (.Y(N171), .A(N135), .B(N134));
NAND2XL inst_cellmath__211__182__I75 (.Y(N172), .A(N141), .B(N140));
INVXL inst_cellmath__211__182__I83 (.Y(N180), .A(N160));
INVXL inst_cellmath__211__182__I84 (.Y(N182), .A(N166));
OAI21XL inst_cellmath__211__182__I85 (.Y(N183), .A0(N165), .A1(N180), .B0(N182));
NOR2XL inst_cellmath__211__182__I87 (.Y(N194), .A(N166), .B(N165));
NAND2BXL inst_cellmath__211__182__I149 (.Y(N189), .AN(N172), .B(N171));
OR2XL inst_cellmath__211__182__I92 (.Y(N191), .A(N172), .B(N171));
OR2XL inst_cellmath__211__182__I97 (.Y(inst_cellmath__211__182__out0[3]), .A(N191), .B(N194));
INVXL inst_cellmath__211__182__I101 (.Y(inst_cellmath__211__182__out0[4]), .A(N191));
OAI21XL inst_cellmath__211__182__I106 (.Y(inst_cellmath__211__182__out0[2]), .A0(N191), .A1(N183), .B0(N189));
AOI21XL inst_cellmath__211__182__I112 (.Y(N216), .A0(N194), .A1(N158), .B0(N164));
OAI2BB1X1 inst_cellmath__211__182__I152 (.Y(N218), .A0N(N140), .A1N(N168), .B0(N141));
OAI21XL inst_cellmath__211__182__I116 (.Y(inst_cellmath__211__182__out0[1]), .A0(N191), .A1(N216), .B0(N218));
OAI21XL inst_cellmath__211__182__I126 (.Y(N232), .A0(N160), .A1(N109), .B0(N115));
OAI21XL inst_cellmath__211__182__I128 (.Y(N234), .A0(N166), .A1(N121), .B0(N127));
AOI21XL inst_cellmath__211__182__I134 (.Y(N240), .A0(N194), .A1(N232), .B0(N234));
OA21X1 inst_cellmath__211__182__I151 (.Y(N242), .A0(N133), .A1(N172), .B0(N139));
OAI21XL inst_cellmath__211__182__I138 (.Y(inst_cellmath__211__182__out0[0]), .A0(N191), .A1(N240), .B0(N242));
endmodule

module cynw_cm_float_cos_inst_cellmath__215_0_bdw1114505291_bdw (
	inst_cellmath__215_0_out0,
	inst_cellmath__215_0_in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__215_0_out0;
input [4:0] inst_cellmath__215_0_in0;
wire N47,N51,N66;
INVXL inst_cellmath__215_0_I64 (.Y(inst_cellmath__215_0_out0[0]), .A(inst_cellmath__215_0_in0[0]));
NAND2XL inst_cellmath__215_0_I21 (.Y(N47), .A(inst_cellmath__215_0_in0[1]), .B(inst_cellmath__215_0_in0[0]));
NAND3XL inst_cellmath__215_0_I23 (.Y(N51), .A(inst_cellmath__215_0_in0[2]), .B(inst_cellmath__215_0_in0[1]), .C(inst_cellmath__215_0_in0[0]));
NAND2BXL inst_cellmath__215_0_I75 (.Y(N66), .AN(inst_cellmath__215_0_in0[3]), .B(N51));
XNOR2X1 inst_cellmath__215_0_I55 (.Y(inst_cellmath__215_0_out0[1]), .A(inst_cellmath__215_0_out0[0]), .B(inst_cellmath__215_0_in0[1]));
XNOR2X1 inst_cellmath__215_0_I56 (.Y(inst_cellmath__215_0_out0[2]), .A(N47), .B(inst_cellmath__215_0_in0[2]));
XOR2XL inst_cellmath__215_0_I76 (.Y(inst_cellmath__215_0_out0[3]), .A(N51), .B(inst_cellmath__215_0_in0[3]));
XNOR2X1 inst_cellmath__215_0_I58 (.Y(inst_cellmath__215_0_out0[4]), .A(N66), .B(inst_cellmath__215_0_in0[4]));
endmodule

module cynw_cm_float_cos_inst_cellmath__220__188__bdw1114505291_bdw (
	inst_cellmath__220__188__out0,
	inst_cellmath__220__188__in0,
	inst_cellmath__220__188__in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__220__188__out0;
input [4:0] inst_cellmath__220__188__in0;
input [47:25] inst_cellmath__220__188__in1;
wire N55,N57,N58,N59,N60,N61,N62 
	,N63,N64,N65,N66,N67,N68,N69,N70 
	,N71,N72,N73,N74,N75,N76,N77,N78 
	,N106,N108,N110,N111,N112,N113,N114,N115 
	,N116,N117,N118,N119,N120,N121,N122,N123 
	,N124,N125,N126,N127,N128,N129,N130,N158 
	,N161,N164,N167,N170,N171,N172,N173,N174 
	,N175,N176,N177,N178,N179,N180,N181,N182 
	,N183,N184,N185,N186,N187,N188,N239,N241 
	,N243,N245,N247,N249,N251,N255,N256,N257 
	,N258,N259,N260,N261,N262,N263,N264,N265 
	,N266,N267,N268,N269,N416,N425,N430,N442 
	,N447,N465,N469,N474,N489;
INVXL inst_cellmath__220__188__I258 (.Y(N416), .A(inst_cellmath__220__188__in0[0]));
AND2XL inst_cellmath__220__188__I2 (.Y(N55), .A(N416), .B(inst_cellmath__220__188__in1[25]));
MX2XL inst_cellmath__220__188__I3 (.Y(N57), .A(inst_cellmath__220__188__in1[25]), .B(inst_cellmath__220__188__in1[26]), .S0(N416));
MX2XL inst_cellmath__220__188__I4 (.Y(N58), .A(inst_cellmath__220__188__in1[26]), .B(inst_cellmath__220__188__in1[27]), .S0(N416));
MX2XL inst_cellmath__220__188__I5 (.Y(N59), .A(inst_cellmath__220__188__in1[27]), .B(inst_cellmath__220__188__in1[28]), .S0(N416));
MX2XL inst_cellmath__220__188__I6 (.Y(N60), .A(inst_cellmath__220__188__in1[28]), .B(inst_cellmath__220__188__in1[29]), .S0(N416));
MX2XL inst_cellmath__220__188__I7 (.Y(N61), .A(inst_cellmath__220__188__in1[29]), .B(inst_cellmath__220__188__in1[30]), .S0(N416));
MX2XL inst_cellmath__220__188__I8 (.Y(N62), .A(inst_cellmath__220__188__in1[30]), .B(inst_cellmath__220__188__in1[31]), .S0(N416));
MX2XL inst_cellmath__220__188__I9 (.Y(N63), .A(inst_cellmath__220__188__in1[31]), .B(inst_cellmath__220__188__in1[32]), .S0(N416));
MX2XL inst_cellmath__220__188__I10 (.Y(N64), .A(inst_cellmath__220__188__in1[32]), .B(inst_cellmath__220__188__in1[33]), .S0(N416));
MX2XL inst_cellmath__220__188__I11 (.Y(N65), .A(inst_cellmath__220__188__in1[33]), .B(inst_cellmath__220__188__in1[34]), .S0(N416));
MX2XL inst_cellmath__220__188__I12 (.Y(N66), .A(inst_cellmath__220__188__in1[34]), .B(inst_cellmath__220__188__in1[35]), .S0(N416));
MX2XL inst_cellmath__220__188__I13 (.Y(N67), .A(inst_cellmath__220__188__in1[35]), .B(inst_cellmath__220__188__in1[36]), .S0(N416));
MX2XL inst_cellmath__220__188__I14 (.Y(N68), .A(inst_cellmath__220__188__in1[36]), .B(inst_cellmath__220__188__in1[37]), .S0(N416));
MX2XL inst_cellmath__220__188__I15 (.Y(N69), .A(inst_cellmath__220__188__in1[37]), .B(inst_cellmath__220__188__in1[38]), .S0(N416));
MX2XL inst_cellmath__220__188__I16 (.Y(N70), .A(inst_cellmath__220__188__in1[38]), .B(inst_cellmath__220__188__in1[39]), .S0(N416));
MX2XL inst_cellmath__220__188__I17 (.Y(N71), .A(inst_cellmath__220__188__in1[39]), .B(inst_cellmath__220__188__in1[40]), .S0(N416));
MX2XL inst_cellmath__220__188__I18 (.Y(N72), .A(inst_cellmath__220__188__in1[40]), .B(inst_cellmath__220__188__in1[41]), .S0(N416));
MX2XL inst_cellmath__220__188__I19 (.Y(N73), .A(inst_cellmath__220__188__in1[41]), .B(inst_cellmath__220__188__in1[42]), .S0(N416));
MX2XL inst_cellmath__220__188__I20 (.Y(N74), .A(inst_cellmath__220__188__in1[42]), .B(inst_cellmath__220__188__in1[43]), .S0(N416));
MX2XL inst_cellmath__220__188__I21 (.Y(N75), .A(inst_cellmath__220__188__in1[43]), .B(inst_cellmath__220__188__in1[44]), .S0(N416));
MX2XL inst_cellmath__220__188__I22 (.Y(N76), .A(inst_cellmath__220__188__in1[44]), .B(inst_cellmath__220__188__in1[45]), .S0(N416));
MX2XL inst_cellmath__220__188__I23 (.Y(N77), .A(inst_cellmath__220__188__in1[45]), .B(inst_cellmath__220__188__in1[46]), .S0(N416));
MX2XL inst_cellmath__220__188__I24 (.Y(N78), .A(inst_cellmath__220__188__in1[46]), .B(inst_cellmath__220__188__in1[47]), .S0(N416));
INVXL inst_cellmath__220__188__I340 (.Y(N425), .A(inst_cellmath__220__188__in0[1]));
INVXL inst_cellmath__220__188__I272 (.Y(N430), .A(N425));
NAND2XL inst_cellmath__220__188__I52 (.Y(N106), .A(N55), .B(N425));
NAND2XL inst_cellmath__220__188__I53 (.Y(N108), .A(N57), .B(N425));
AOI22XL inst_cellmath__220__188__I54 (.Y(N110), .A0(N430), .A1(N55), .B0(N58), .B1(N425));
AOI22XL inst_cellmath__220__188__I55 (.Y(N111), .A0(N430), .A1(N57), .B0(N59), .B1(N425));
AOI22XL inst_cellmath__220__188__I56 (.Y(N112), .A0(N430), .A1(N58), .B0(N60), .B1(N425));
AOI22XL inst_cellmath__220__188__I57 (.Y(N113), .A0(N430), .A1(N59), .B0(N61), .B1(N425));
AOI22XL inst_cellmath__220__188__I58 (.Y(N114), .A0(N430), .A1(N60), .B0(N62), .B1(N425));
AOI22XL inst_cellmath__220__188__I59 (.Y(N115), .A0(N430), .A1(N61), .B0(N63), .B1(N425));
AOI22XL inst_cellmath__220__188__I60 (.Y(N116), .A0(N430), .A1(N62), .B0(N64), .B1(N425));
AOI22XL inst_cellmath__220__188__I61 (.Y(N117), .A0(N430), .A1(N63), .B0(N65), .B1(N425));
AOI22XL inst_cellmath__220__188__I62 (.Y(N118), .A0(N430), .A1(N64), .B0(N66), .B1(N425));
AOI22XL inst_cellmath__220__188__I63 (.Y(N119), .A0(N430), .A1(N65), .B0(N67), .B1(N425));
AOI22XL inst_cellmath__220__188__I64 (.Y(N120), .A0(N430), .A1(N66), .B0(N68), .B1(N425));
AOI22XL inst_cellmath__220__188__I65 (.Y(N121), .A0(N430), .A1(N67), .B0(N69), .B1(N425));
AOI22XL inst_cellmath__220__188__I66 (.Y(N122), .A0(N430), .A1(N68), .B0(N70), .B1(N425));
AOI22XL inst_cellmath__220__188__I67 (.Y(N123), .A0(N430), .A1(N69), .B0(N71), .B1(N425));
AOI22XL inst_cellmath__220__188__I68 (.Y(N124), .A0(N430), .A1(N70), .B0(N72), .B1(N425));
AOI22XL inst_cellmath__220__188__I69 (.Y(N125), .A0(N430), .A1(N71), .B0(N73), .B1(N425));
AOI22XL inst_cellmath__220__188__I70 (.Y(N126), .A0(N430), .A1(N72), .B0(N74), .B1(N425));
AOI22XL inst_cellmath__220__188__I71 (.Y(N127), .A0(N430), .A1(N73), .B0(N75), .B1(N425));
AOI22XL inst_cellmath__220__188__I72 (.Y(N128), .A0(N430), .A1(N74), .B0(N76), .B1(N425));
AOI22XL inst_cellmath__220__188__I73 (.Y(N129), .A0(N430), .A1(N75), .B0(N77), .B1(N425));
AOI22XL inst_cellmath__220__188__I74 (.Y(N130), .A0(N430), .A1(N76), .B0(N78), .B1(N425));
INVXL inst_cellmath__220__188__I341 (.Y(N442), .A(inst_cellmath__220__188__in0[2]));
INVXL inst_cellmath__220__188__I289 (.Y(N447), .A(N442));
NOR2XL inst_cellmath__220__188__I102 (.Y(N158), .A(N447), .B(N106));
NOR2XL inst_cellmath__220__188__I103 (.Y(N161), .A(N447), .B(N108));
NOR2XL inst_cellmath__220__188__I104 (.Y(N164), .A(N447), .B(N110));
NOR2XL inst_cellmath__220__188__I105 (.Y(N167), .A(N447), .B(N111));
AOI22XL inst_cellmath__220__188__I106 (.Y(N170), .A0(N442), .A1(N112), .B0(N106), .B1(N447));
AOI22XL inst_cellmath__220__188__I107 (.Y(N171), .A0(N442), .A1(N113), .B0(N108), .B1(N447));
AOI22XL inst_cellmath__220__188__I108 (.Y(N172), .A0(N442), .A1(N114), .B0(N110), .B1(N447));
AOI22XL inst_cellmath__220__188__I109 (.Y(N173), .A0(N442), .A1(N115), .B0(N111), .B1(N447));
AOI22XL inst_cellmath__220__188__I110 (.Y(N174), .A0(N442), .A1(N116), .B0(N112), .B1(N447));
AOI22XL inst_cellmath__220__188__I111 (.Y(N175), .A0(N442), .A1(N117), .B0(N113), .B1(N447));
AOI22XL inst_cellmath__220__188__I112 (.Y(N176), .A0(N442), .A1(N118), .B0(N114), .B1(N447));
AOI22XL inst_cellmath__220__188__I113 (.Y(N177), .A0(N442), .A1(N119), .B0(N115), .B1(N447));
AOI22XL inst_cellmath__220__188__I114 (.Y(N178), .A0(N442), .A1(N120), .B0(N116), .B1(N447));
AOI22XL inst_cellmath__220__188__I115 (.Y(N179), .A0(N442), .A1(N121), .B0(N117), .B1(N447));
AOI22XL inst_cellmath__220__188__I116 (.Y(N180), .A0(N442), .A1(N122), .B0(N118), .B1(N447));
AOI22XL inst_cellmath__220__188__I117 (.Y(N181), .A0(N442), .A1(N123), .B0(N119), .B1(N447));
AOI22XL inst_cellmath__220__188__I118 (.Y(N182), .A0(N442), .A1(N124), .B0(N120), .B1(N447));
AOI22XL inst_cellmath__220__188__I119 (.Y(N183), .A0(N442), .A1(N125), .B0(N121), .B1(N447));
AOI22XL inst_cellmath__220__188__I120 (.Y(N184), .A0(N442), .A1(N126), .B0(N122), .B1(N447));
AOI22XL inst_cellmath__220__188__I121 (.Y(N185), .A0(N442), .A1(N127), .B0(N123), .B1(N447));
AOI22XL inst_cellmath__220__188__I122 (.Y(N186), .A0(N442), .A1(N128), .B0(N124), .B1(N447));
AOI22XL inst_cellmath__220__188__I123 (.Y(N187), .A0(N442), .A1(N129), .B0(N125), .B1(N447));
AOI22XL inst_cellmath__220__188__I124 (.Y(N188), .A0(N442), .A1(N130), .B0(N126), .B1(N447));
INVXL inst_cellmath__220__188__I307 (.Y(N465), .A(inst_cellmath__220__188__in0[3]));
NAND2XL inst_cellmath__220__188__I152 (.Y(N239), .A(N158), .B(N465));
NAND2XL inst_cellmath__220__188__I153 (.Y(N241), .A(N161), .B(N465));
NAND2XL inst_cellmath__220__188__I154 (.Y(N243), .A(N164), .B(N465));
NAND2XL inst_cellmath__220__188__I155 (.Y(N245), .A(N167), .B(N465));
NAND2XL inst_cellmath__220__188__I156 (.Y(N247), .A(N170), .B(N465));
NAND2XL inst_cellmath__220__188__I157 (.Y(N249), .A(N171), .B(N465));
NAND2XL inst_cellmath__220__188__I158 (.Y(N251), .A(N172), .B(N465));
AOI22XL inst_cellmath__220__188__I160 (.Y(N255), .A0(inst_cellmath__220__188__in0[3]), .A1(N158), .B0(N174), .B1(N465));
AOI22XL inst_cellmath__220__188__I161 (.Y(N256), .A0(inst_cellmath__220__188__in0[3]), .A1(N161), .B0(N175), .B1(N465));
AOI22XL inst_cellmath__220__188__I162 (.Y(N257), .A0(inst_cellmath__220__188__in0[3]), .A1(N164), .B0(N176), .B1(N465));
AOI22XL inst_cellmath__220__188__I163 (.Y(N258), .A0(inst_cellmath__220__188__in0[3]), .A1(N167), .B0(N177), .B1(N465));
AOI22XL inst_cellmath__220__188__I164 (.Y(N259), .A0(inst_cellmath__220__188__in0[3]), .A1(N170), .B0(N178), .B1(N465));
AOI22XL inst_cellmath__220__188__I165 (.Y(N260), .A0(inst_cellmath__220__188__in0[3]), .A1(N171), .B0(N179), .B1(N465));
AOI22XL inst_cellmath__220__188__I166 (.Y(N261), .A0(inst_cellmath__220__188__in0[3]), .A1(N172), .B0(N180), .B1(N465));
AOI22XL inst_cellmath__220__188__I167 (.Y(N262), .A0(inst_cellmath__220__188__in0[3]), .A1(N173), .B0(N181), .B1(N465));
AOI22XL inst_cellmath__220__188__I168 (.Y(N263), .A0(inst_cellmath__220__188__in0[3]), .A1(N174), .B0(N182), .B1(N465));
AOI22XL inst_cellmath__220__188__I169 (.Y(N264), .A0(inst_cellmath__220__188__in0[3]), .A1(N175), .B0(N183), .B1(N465));
AOI22XL inst_cellmath__220__188__I170 (.Y(N265), .A0(inst_cellmath__220__188__in0[3]), .A1(N176), .B0(N184), .B1(N465));
AOI22XL inst_cellmath__220__188__I171 (.Y(N266), .A0(inst_cellmath__220__188__in0[3]), .A1(N177), .B0(N185), .B1(N465));
AOI22XL inst_cellmath__220__188__I172 (.Y(N267), .A0(inst_cellmath__220__188__in0[3]), .A1(N178), .B0(N186), .B1(N465));
AOI22XL inst_cellmath__220__188__I173 (.Y(N268), .A0(inst_cellmath__220__188__in0[3]), .A1(N179), .B0(N187), .B1(N465));
AOI22XL inst_cellmath__220__188__I174 (.Y(N269), .A0(inst_cellmath__220__188__in0[3]), .A1(N180), .B0(N188), .B1(N465));
INVXL inst_cellmath__220__188__I337 (.Y(N469), .A(inst_cellmath__220__188__in0[4]));
INVXL inst_cellmath__220__188__I316 (.Y(N474), .A(N469));
NOR2XL inst_cellmath__220__188__I202 (.Y(inst_cellmath__220__188__out0[0]), .A(N474), .B(N239));
NOR2XL inst_cellmath__220__188__I203 (.Y(inst_cellmath__220__188__out0[1]), .A(N474), .B(N241));
NOR2XL inst_cellmath__220__188__I204 (.Y(inst_cellmath__220__188__out0[2]), .A(N474), .B(N243));
NOR2XL inst_cellmath__220__188__I205 (.Y(inst_cellmath__220__188__out0[3]), .A(N474), .B(N245));
NOR2XL inst_cellmath__220__188__I206 (.Y(inst_cellmath__220__188__out0[4]), .A(N474), .B(N247));
NOR2XL inst_cellmath__220__188__I207 (.Y(inst_cellmath__220__188__out0[5]), .A(N474), .B(N249));
NOR2XL inst_cellmath__220__188__I208 (.Y(inst_cellmath__220__188__out0[6]), .A(N474), .B(N251));
NAND2XL hyperpropagate_3_1_A_I342 (.Y(N489), .A(N173), .B(N465));
NOR2XL hyperpropagate_3_1_A_I343 (.Y(inst_cellmath__220__188__out0[7]), .A(N474), .B(N489));
NOR2XL inst_cellmath__220__188__I210 (.Y(inst_cellmath__220__188__out0[8]), .A(N474), .B(N255));
NOR2XL inst_cellmath__220__188__I211 (.Y(inst_cellmath__220__188__out0[9]), .A(N474), .B(N256));
NOR2XL inst_cellmath__220__188__I212 (.Y(inst_cellmath__220__188__out0[10]), .A(N474), .B(N257));
NOR2XL inst_cellmath__220__188__I213 (.Y(inst_cellmath__220__188__out0[11]), .A(N474), .B(N258));
NOR2XL inst_cellmath__220__188__I214 (.Y(inst_cellmath__220__188__out0[12]), .A(N474), .B(N259));
NOR2XL inst_cellmath__220__188__I215 (.Y(inst_cellmath__220__188__out0[13]), .A(N474), .B(N260));
NOR2XL inst_cellmath__220__188__I216 (.Y(inst_cellmath__220__188__out0[14]), .A(N474), .B(N261));
NOR2XL inst_cellmath__220__188__I217 (.Y(inst_cellmath__220__188__out0[15]), .A(N474), .B(N262));
AOI22XL inst_cellmath__220__188__I218 (.Y(inst_cellmath__220__188__out0[16]), .A0(N469), .A1(N263), .B0(N239), .B1(N474));
AOI22XL inst_cellmath__220__188__I219 (.Y(inst_cellmath__220__188__out0[17]), .A0(N469), .A1(N264), .B0(N241), .B1(N474));
AOI22XL inst_cellmath__220__188__I220 (.Y(inst_cellmath__220__188__out0[18]), .A0(N469), .A1(N265), .B0(N243), .B1(N474));
AOI22XL inst_cellmath__220__188__I221 (.Y(inst_cellmath__220__188__out0[19]), .A0(N469), .A1(N266), .B0(N245), .B1(N474));
AOI22XL inst_cellmath__220__188__I222 (.Y(inst_cellmath__220__188__out0[20]), .A0(N469), .A1(N267), .B0(N247), .B1(N474));
AOI22XL inst_cellmath__220__188__I223 (.Y(inst_cellmath__220__188__out0[21]), .A0(N469), .A1(N268), .B0(N249), .B1(N474));
AOI22XL inst_cellmath__220__188__I224 (.Y(inst_cellmath__220__188__out0[22]), .A0(N469), .A1(N269), .B0(N251), .B1(N474));
endmodule

module cynw_cm_float_cos_inst_cellmath__221__195__bdw1114505291_bdw (
	inst_cellmath__221__195__out0,
	inst_cellmath__221__195__in0
	); /* architecture "gate_level" */ 
output [6:0] inst_cellmath__221__195__out0;
input [4:0] inst_cellmath__221__195__in0;
INVXL inst_cellmath__221__195__I5 (.Y(inst_cellmath__221__195__out0[0]), .A(inst_cellmath__221__195__in0[0]));
INVXL inst_cellmath__221__195__I6 (.Y(inst_cellmath__221__195__out0[1]), .A(inst_cellmath__221__195__in0[1]));
INVXL inst_cellmath__221__195__I7 (.Y(inst_cellmath__221__195__out0[2]), .A(inst_cellmath__221__195__in0[2]));
INVXL inst_cellmath__221__195__I8 (.Y(inst_cellmath__221__195__out0[3]), .A(inst_cellmath__221__195__in0[3]));
INVXL inst_cellmath__221__195__I9 (.Y(inst_cellmath__221__195__out0[4]), .A(inst_cellmath__221__195__in0[4]));
assign inst_cellmath__221__195__out0[5] = 1'B1;
assign inst_cellmath__221__195__out0[6] = 1'B1;
endmodule

module cynw_cm_float_cos_inst_cellmath__220_2WWMM_bdw1114505291_bdw (
	inst_cellmath__220_2WWMM_out0,
	inst_cellmath__220_2WWMM_in0,
	inst_cellmath__220_2WWMM_in1,
	inst_cellmath__220_2WWMM_in2
	); /* architecture "gate_level" */ 
output [30:0] inst_cellmath__220_2WWMM_out0;
input [6:0] inst_cellmath__220_2WWMM_in0;
input [22:0] inst_cellmath__220_2WWMM_in1;
input  inst_cellmath__220_2WWMM_in2;
wire N168;
INVXL inst_cellmath__220_2WWMM_I34 (.Y(N168), .A(inst_cellmath__220_2WWMM_in2));
NAND2BXL inst_cellmath__220_2WWMM_I1 (.Y(inst_cellmath__220_2WWMM_out0[0]), .AN(inst_cellmath__220_2WWMM_in0[0]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I2 (.Y(inst_cellmath__220_2WWMM_out0[1]), .AN(inst_cellmath__220_2WWMM_in0[1]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I3 (.Y(inst_cellmath__220_2WWMM_out0[2]), .AN(inst_cellmath__220_2WWMM_in0[2]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I4 (.Y(inst_cellmath__220_2WWMM_out0[3]), .AN(inst_cellmath__220_2WWMM_in0[3]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I5 (.Y(inst_cellmath__220_2WWMM_out0[4]), .AN(inst_cellmath__220_2WWMM_in0[4]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I6 (.Y(inst_cellmath__220_2WWMM_out0[5]), .AN(inst_cellmath__220_2WWMM_in0[5]), .B(N168));
NAND2BXL inst_cellmath__220_2WWMM_I7 (.Y(inst_cellmath__220_2WWMM_out0[6]), .AN(inst_cellmath__220_2WWMM_in0[6]), .B(N168));
AND2XL inst_cellmath__220_2WWMM_I9 (.Y(inst_cellmath__220_2WWMM_out0[8]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[0]));
AND2XL inst_cellmath__220_2WWMM_I10 (.Y(inst_cellmath__220_2WWMM_out0[9]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[1]));
AND2XL inst_cellmath__220_2WWMM_I11 (.Y(inst_cellmath__220_2WWMM_out0[10]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[2]));
AND2XL inst_cellmath__220_2WWMM_I12 (.Y(inst_cellmath__220_2WWMM_out0[11]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[3]));
AND2XL inst_cellmath__220_2WWMM_I13 (.Y(inst_cellmath__220_2WWMM_out0[12]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[4]));
AND2XL inst_cellmath__220_2WWMM_I14 (.Y(inst_cellmath__220_2WWMM_out0[13]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[5]));
AND2XL inst_cellmath__220_2WWMM_I15 (.Y(inst_cellmath__220_2WWMM_out0[14]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[6]));
AND2XL inst_cellmath__220_2WWMM_I16 (.Y(inst_cellmath__220_2WWMM_out0[15]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[7]));
AND2XL inst_cellmath__220_2WWMM_I17 (.Y(inst_cellmath__220_2WWMM_out0[16]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[8]));
AND2XL inst_cellmath__220_2WWMM_I18 (.Y(inst_cellmath__220_2WWMM_out0[17]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[9]));
AND2XL inst_cellmath__220_2WWMM_I19 (.Y(inst_cellmath__220_2WWMM_out0[18]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[10]));
AND2XL inst_cellmath__220_2WWMM_I20 (.Y(inst_cellmath__220_2WWMM_out0[19]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[11]));
AND2XL inst_cellmath__220_2WWMM_I21 (.Y(inst_cellmath__220_2WWMM_out0[20]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[12]));
AND2XL inst_cellmath__220_2WWMM_I22 (.Y(inst_cellmath__220_2WWMM_out0[21]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[13]));
AND2XL inst_cellmath__220_2WWMM_I23 (.Y(inst_cellmath__220_2WWMM_out0[22]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[14]));
AND2XL inst_cellmath__220_2WWMM_I24 (.Y(inst_cellmath__220_2WWMM_out0[23]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[15]));
AND2XL inst_cellmath__220_2WWMM_I25 (.Y(inst_cellmath__220_2WWMM_out0[24]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[16]));
AND2XL inst_cellmath__220_2WWMM_I26 (.Y(inst_cellmath__220_2WWMM_out0[25]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[17]));
AND2XL inst_cellmath__220_2WWMM_I27 (.Y(inst_cellmath__220_2WWMM_out0[26]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[18]));
AND2XL inst_cellmath__220_2WWMM_I28 (.Y(inst_cellmath__220_2WWMM_out0[27]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[19]));
AND2XL inst_cellmath__220_2WWMM_I29 (.Y(inst_cellmath__220_2WWMM_out0[28]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[20]));
AND2XL inst_cellmath__220_2WWMM_I30 (.Y(inst_cellmath__220_2WWMM_out0[29]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[21]));
AND2XL inst_cellmath__220_2WWMM_I31 (.Y(inst_cellmath__220_2WWMM_out0[30]), .A(N168), .B(inst_cellmath__220_2WWMM_in1[22]));
assign inst_cellmath__220_2WWMM_out0[7] = 1'B0;
endmodule

module cynw_cm_float_cos_inst_cellmath__223__208__bdw1114505291_bdw (
	inst_cellmath__223__208__out0,
	inst_cellmath__223__208__in0,
	inst_cellmath__223__208__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__208__out0;
input [6:0] inst_cellmath__223__208__in0;
input [29:8] inst_cellmath__223__208__in1;
wire N37,N38,N39,N41,N46,N47,N48 
	,N50,N51,N53,N59,N61,N64,N65,N67 
	;
OR4X1 inst_cellmath__223__208__I40 (.Y(N37), .A(inst_cellmath__223__208__in0[6]), .B(inst_cellmath__223__208__in0[5]), .C(inst_cellmath__223__208__in0[0]), .D(inst_cellmath__223__208__in0[1]));
NOR2XL inst_cellmath__223__208__I6 (.Y(N38), .A(N37), .B(inst_cellmath__223__208__in0[2]));
NOR2XL inst_cellmath__223__208__I7 (.Y(N39), .A(inst_cellmath__223__208__in0[3]), .B(inst_cellmath__223__208__in0[4]));
NAND3BXL inst_cellmath__223__208__I41 (.Y(N41), .AN(inst_cellmath__223__208__in1[9]), .B(N39), .C(N38));
OR4X1 inst_cellmath__223__208__I43 (.Y(N46), .A(inst_cellmath__223__208__in1[8]), .B(inst_cellmath__223__208__in1[10]), .C(N41), .D(inst_cellmath__223__208__in1[11]));
NOR2XL inst_cellmath__223__208__I15 (.Y(N47), .A(inst_cellmath__223__208__in1[15]), .B(inst_cellmath__223__208__in1[12]));
NOR2XL inst_cellmath__223__208__I16 (.Y(N48), .A(inst_cellmath__223__208__in1[14]), .B(inst_cellmath__223__208__in1[13]));
NOR2XL inst_cellmath__223__208__I18 (.Y(N50), .A(inst_cellmath__223__208__in1[16]), .B(inst_cellmath__223__208__in1[18]));
NOR2XL inst_cellmath__223__208__I19 (.Y(N51), .A(inst_cellmath__223__208__in1[17]), .B(inst_cellmath__223__208__in1[23]));
NAND2XL inst_cellmath__223__208__I21 (.Y(N53), .A(N47), .B(N48));
NOR3XL inst_cellmath__223__208__I44 (.Y(N65), .A(inst_cellmath__223__208__in1[20]), .B(inst_cellmath__223__208__in1[19]), .C(inst_cellmath__223__208__in1[28]));
NAND2XL inst_cellmath__223__208__I27 (.Y(N59), .A(N50), .B(N51));
NOR3XL inst_cellmath__223__208__I45 (.Y(N61), .A(inst_cellmath__223__208__in1[22]), .B(inst_cellmath__223__208__in1[21]), .C(N53));
NOR4X1 inst_cellmath__223__208__I50 (.Y(N67), .A(inst_cellmath__223__208__in1[25]), .B(inst_cellmath__223__208__in1[27]), .C(inst_cellmath__223__208__in1[29]), .D(N46));
NOR3XL inst_cellmath__223__208__I47 (.Y(N64), .A(inst_cellmath__223__208__in1[24]), .B(inst_cellmath__223__208__in1[26]), .C(N59));
NAND4XL inst_cellmath__223__208__I92 (.Y(inst_cellmath__223__208__out0[0]), .A(N64), .B(N61), .C(N65), .D(N67));
endmodule

module cynw_cm_float_cos_inst_cellmath__223__199__bdw1114505291_bdw (
	inst_cellmath__223__199__out0,
	inst_cellmath__223__199__in0,
	inst_cellmath__223__199__in1,
	inst_cellmath__223__199__in2,
	inst_cellmath__223__199__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__199__out0;
input  inst_cellmath__223__199__in0;
input [1:1] inst_cellmath__223__199__in1;
input [8:6] inst_cellmath__223__199__in2;
input [0:0] inst_cellmath__223__199__in3;
wire N9,N10;
NOR2XL inst_cellmath__223__199__I0 (.Y(N9), .A(inst_cellmath__223__199__in2[8]), .B(inst_cellmath__223__199__in2[7]));
NOR2XL inst_cellmath__223__199__I1 (.Y(N10), .A(inst_cellmath__223__199__in2[6]), .B(inst_cellmath__223__199__in0));
AND4XL inst_cellmath__223__199__I16 (.Y(inst_cellmath__223__199__out0[0]), .A(N9), .B(N10), .C(inst_cellmath__223__199__in1[1]), .D(inst_cellmath__223__199__in3[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__224__213__bdw1114505291_bdw (
	inst_cellmath__224__213__out0,
	inst_cellmath__224__213__in0,
	inst_cellmath__224__213__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__224__213__out0;
input [0:0] inst_cellmath__224__213__in0;
input  inst_cellmath__224__213__in1;
OR2XL inst_cellmath__224__213__I0 (.Y(inst_cellmath__224__213__out0[0]), .A(inst_cellmath__224__213__in1), .B(inst_cellmath__224__213__in0[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__224__212__bdw1114505291_bdw (
	inst_cellmath__224__212__out0,
	inst_cellmath__224__212__in0,
	inst_cellmath__224__212__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__224__212__out0;
input  inst_cellmath__224__212__in0;
input [0:0] inst_cellmath__224__212__in1;
NAND2BXL inst_cellmath__224__212__I2 (.Y(inst_cellmath__224__212__out0[0]), .AN(inst_cellmath__224__212__in0), .B(inst_cellmath__224__212__in1[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__225__215__bdw1114505291_bdw (
	inst_cellmath__225__215__out0,
	inst_cellmath__225__215__in0,
	inst_cellmath__225__215__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__225__215__out0;
input  inst_cellmath__225__215__in0,
	inst_cellmath__225__215__in1;
NAND2BXL inst_cellmath__225__215__I2 (.Y(inst_cellmath__225__215__out0[0]), .AN(inst_cellmath__225__215__in0), .B(inst_cellmath__225__215__in1));
endmodule

module cynw_cm_float_cos_inst_cellmath__228_0_bdw1114505291_bdw (
	inst_cellmath__228_0_out0,
	inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1,
	inst_cellmath__228_0_in2,
	inst_cellmath__228_0_in3
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__228_0_out0;
input [0:0] inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1,
	inst_cellmath__228_0_in2;
input [6:0] inst_cellmath__228_0_in3;
wire N92,N100;
INVXL buf1_A_I40 (.Y(N100), .A(inst_cellmath__228_0_in0[0]));
INVXL buf1_A_I41 (.Y(N92), .A(N100));
MX2XL inst_cellmath__228_0_I16 (.Y(inst_cellmath__228_0_out0[0]), .A(inst_cellmath__228_0_in3[0]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I17 (.Y(inst_cellmath__228_0_out0[1]), .A(inst_cellmath__228_0_in3[1]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I18 (.Y(inst_cellmath__228_0_out0[2]), .A(inst_cellmath__228_0_in3[2]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I19 (.Y(inst_cellmath__228_0_out0[3]), .A(inst_cellmath__228_0_in3[3]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I20 (.Y(inst_cellmath__228_0_out0[4]), .A(inst_cellmath__228_0_in3[4]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I21 (.Y(inst_cellmath__228_0_out0[5]), .A(inst_cellmath__228_0_in3[5]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
MX2XL inst_cellmath__228_0_I22 (.Y(inst_cellmath__228_0_out0[6]), .A(inst_cellmath__228_0_in3[6]), .B(inst_cellmath__228_0_in1[0]), .S0(N92));
AND2XL inst_cellmath__228_0_I36 (.Y(inst_cellmath__228_0_out0[7]), .A(N92), .B(inst_cellmath__228_0_in2[0]));
endmodule

module cynw_cm_float_cos_inst_cellmath__231_0_bdw1114505291_bdw (
	inst_cellmath__231_0_out0,
	inst_cellmath__231_0_in0,
	inst_cellmath__231_0_in1,
	inst_cellmath__231_0_in2,
	inst_cellmath__231_0_in3
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__231_0_out0;
input  inst_cellmath__231_0_in0;
input [0:0] inst_cellmath__231_0_in1;
input [30:8] inst_cellmath__231_0_in2;
input [46:46] inst_cellmath__231_0_in3;
MX2XL inst_cellmath__231_0_I46 (.Y(inst_cellmath__231_0_out0[0]), .A(inst_cellmath__231_0_in2[8]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I47 (.Y(inst_cellmath__231_0_out0[1]), .A(inst_cellmath__231_0_in2[9]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I48 (.Y(inst_cellmath__231_0_out0[2]), .A(inst_cellmath__231_0_in2[10]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I49 (.Y(inst_cellmath__231_0_out0[3]), .A(inst_cellmath__231_0_in2[11]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I50 (.Y(inst_cellmath__231_0_out0[4]), .A(inst_cellmath__231_0_in2[12]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I51 (.Y(inst_cellmath__231_0_out0[5]), .A(inst_cellmath__231_0_in2[13]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I52 (.Y(inst_cellmath__231_0_out0[6]), .A(inst_cellmath__231_0_in2[14]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I53 (.Y(inst_cellmath__231_0_out0[7]), .A(inst_cellmath__231_0_in2[15]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I54 (.Y(inst_cellmath__231_0_out0[8]), .A(inst_cellmath__231_0_in2[16]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I55 (.Y(inst_cellmath__231_0_out0[9]), .A(inst_cellmath__231_0_in2[17]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I56 (.Y(inst_cellmath__231_0_out0[10]), .A(inst_cellmath__231_0_in2[18]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I57 (.Y(inst_cellmath__231_0_out0[11]), .A(inst_cellmath__231_0_in2[19]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I58 (.Y(inst_cellmath__231_0_out0[12]), .A(inst_cellmath__231_0_in2[20]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I59 (.Y(inst_cellmath__231_0_out0[13]), .A(inst_cellmath__231_0_in2[21]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I60 (.Y(inst_cellmath__231_0_out0[14]), .A(inst_cellmath__231_0_in2[22]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I61 (.Y(inst_cellmath__231_0_out0[15]), .A(inst_cellmath__231_0_in2[23]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I62 (.Y(inst_cellmath__231_0_out0[16]), .A(inst_cellmath__231_0_in2[24]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I63 (.Y(inst_cellmath__231_0_out0[17]), .A(inst_cellmath__231_0_in2[25]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I64 (.Y(inst_cellmath__231_0_out0[18]), .A(inst_cellmath__231_0_in2[26]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I65 (.Y(inst_cellmath__231_0_out0[19]), .A(inst_cellmath__231_0_in2[27]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I66 (.Y(inst_cellmath__231_0_out0[20]), .A(inst_cellmath__231_0_in2[28]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I67 (.Y(inst_cellmath__231_0_out0[21]), .A(inst_cellmath__231_0_in2[29]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
MX2XL inst_cellmath__231_0_I68 (.Y(inst_cellmath__231_0_out0[22]), .A(inst_cellmath__231_0_in2[30]), .B(inst_cellmath__231_0_in0), .S0(inst_cellmath__231_0_in1[0]));
endmodule

/* CADENCE  vrH0TAjfrBk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




module DFT_compute_cynw_cm_float_cos_E8_M23_4( a_sign, a_exp, a_man, x, aclk, astall );
input a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire[36:0] x_wire;
input aclk;
input astall;
cynw_cm_float_cos_inst_cellmath__231_0_bdw1114505291_bdw cynw_cm_float_cos_inst_cellmath__231_0_bdw2869798270_bdw_inst( .a_sign(a_sign), .a_exp(a_exp), .a_man(a_man), .x(x_wire));
reg [36:0] x_reg_0;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_0 <= x_wire;
end
/* $A : movable_reg = reset */
reg [36:0] x_reg_1;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_1 <= x_reg_0;
end
/* $A : movable_reg = reset */
assign x = x_reg_1;
endmodule


