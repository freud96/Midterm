/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:43 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_add2_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40;
wire [8:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49;
wire [25:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52;
wire [5:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55;
wire [25:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62;
wire [24:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63;
wire [7:0] DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66;
wire  DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417,
	DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423;
wire N3881,N4038,N4247,N4249,N4293,N4572,N4578 
	,N4892,N4894,N4901,N4903,N5139,N5145,N5154,N5398 
	,N5409,N5467,N5475,N5508,N5977,N5979,N5981,N5984 
	,N5986,N5988,N6007,N6009,N6073,N6075,N6077,N6083 
	,N6087,N6089,N6097,N6101,N6107,N6109,N6113,N6122 
	,N6124,N6129,N6133,N6135,N6143,N6147,N6156,N6158 
	,N6173,N6175,N6185,N6192,N6194,N6201,N6203,N6210 
	,N6212,N6217,N6221,N6228,N6230,N6235,N6239,N6246 
	,N6248,N6253,N6257,N6262,N6266,N6271,N6275,N6280 
	,N6284,N6289,N6295,N6298,N6304,N6331,N6341,N6349 
	,N6355,N6364,N6370,N6654,N6657,N6663,N6666,N6675 
	,N6677,N6853,N6854,N6856,N6863,N6870,N6918;
EDFFHQX1 x_reg_23__retimed_I3276 (.Q(N6677), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3275 (.Q(N6675), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_29__retimed_I3271 (.Q(N6666), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_27__retimed_I3270 (.Q(N6663), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3268 (.Q(N6657), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I3267 (.Q(N6654), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3144 (.Q(N6304), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3141 (.Q(N6298), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3140 (.Q(N6295), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3137 (.Q(N6289), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3135 (.Q(N6284), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3133 (.Q(N6280), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3131 (.Q(N6275), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3129 (.Q(N6271), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3127 (.Q(N6266), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3125 (.Q(N6262), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3123 (.Q(N6257), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3121 (.Q(N6253), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3119 (.Q(N6248), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3118 (.Q(N6246), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3115 (.Q(N6239), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3113 (.Q(N6235), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3111 (.Q(N6230), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3110 (.Q(N6228), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3107 (.Q(N6221), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3105 (.Q(N6217), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3103 (.Q(N6212), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3102 (.Q(N6210), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3099 (.Q(N6203), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3098 (.Q(N6201), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3095 (.Q(N6194), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3094 (.Q(N6192), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3091 (.Q(N6185), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3089 (.Q(N6175), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3088 (.Q(N6173), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3084 (.Q(N6158), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3083 (.Q(N6156), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3080 (.Q(N6147), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3078 (.Q(N6143), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3076 (.Q(N6135), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3075 (.Q(N6133), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3073 (.Q(N6129), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3072 (.Q(N6124), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3071 (.Q(N6122), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3068 (.Q(N6113), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3066 (.Q(N6109), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3065 (.Q(N6107), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3064 (.Q(N6101), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3062 (.Q(N6097), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3060 (.Q(N6089), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3059 (.Q(N6087), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3057 (.Q(N6083), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3056 (.Q(N6077), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3055 (.Q(N6075), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435), .E(bdw_enable), .CK(aclk));
EDFFHQX2 x_reg_30__retimed_I3054 (.Q(N6073), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3041 (.Q(N6009), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I3040 (.Q(N6007), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3036 (.Q(N5988), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3035 (.Q(N5986), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420), .E(bdw_enable), .CK(aclk));
EDFFHQX2 x_reg_23__retimed_I3034 (.Q(N5984), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3033 (.Q(N5981), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3032 (.Q(N5979), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I3031 (.Q(N5977), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I2872 (.Q(N5508), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I2861 (.Q(N5475), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2858 (.Q(N5467), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2849 (.Q(N5409), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_25__retimed_I2844 (.Q(N5398), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2767 (.Q(N5154), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_26__retimed_I2763 (.Q(N5145), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2761 (.Q(N5139), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I2682 (.Q(N4903), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I2681 (.Q(N4901), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2678 (.Q(N4894), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2677 (.Q(N4892), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_28__retimed_I2572 (.Q(N4578), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2570 (.Q(N4572), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2465 (.Q(N4293), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I2460 (.Q(N4249), .D(b_sign), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_31__retimed_I2459 (.Q(N4247), .D(a_sign), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_30__retimed_I2367 (.Q(N4038), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I2300 (.Q(N3881), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62), .E(bdw_enable), .CK(aclk));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3363 (.Y(N6853), .A(N3881));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3364 (.Y(N6854), .A(N6853));
INVX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I0 (.Y(bdw_enable), .A(astall));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I1 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131), .A(b_exp[0]), .B(b_exp[1]));
AND4XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I2 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187), .A(b_exp[7]), .B(b_exp[6]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3133));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I4 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3131), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6187));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I5 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I6 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3167));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I7 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154), .A(b_man[10]), .B(b_man[9]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I8 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173), .A(b_man[6]), .B(b_man[5]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I9 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162), .A(b_man[8]), .B(b_man[7]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I10 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182), .A(b_man[4]), .B(b_man[3]));
NAND4XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I11 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3154), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3173), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3162), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3182));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I12 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I13 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I14 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3171), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3165), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3176), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3186));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I15 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I16 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018), .A(a_exp[0]));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I17 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10018));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I18 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019), .B(a_exp[1]));
AND4XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I19 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I20 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195), .A(a_exp[7]), .B(a_exp[6]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3222));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I21 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3220), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6195));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I22 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I23 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3256));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I24 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243), .A(a_man[10]), .B(a_man[9]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I25 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262), .A(a_man[6]), .B(a_man[5]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I26 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251), .A(a_man[8]), .B(a_man[7]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I27 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271), .A(a_man[4]), .B(a_man[3]));
NAND4XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I28 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3243), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3262), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3251), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3271));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I29 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I30 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I31 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3260), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3254), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3265), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3275));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I32 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I33 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__30), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__32));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I34 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__27), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__29));
XOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I35 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .A(a_sign), .B(b_sign));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I36 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__24), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__21), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]));
OR3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I37 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__62), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__23), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__20), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N495));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I38 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I39 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I40 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I41 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3010), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3014));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I42 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988), .A(a_exp[7]), .B(a_exp[1]), .C(a_exp[6]), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I43 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I44 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2988), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2992));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I45 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I46 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504), .A(a_exp[4]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I47 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362), .A(a_exp[3]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I48 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502), .A(a_exp[2]));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I49 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501), .A(a_exp[1]));
INVX2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I50 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500), .A(a_exp[0]));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I51 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178), .A(b_exp[0]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I52 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6178));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I53 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[1]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501), .B(b_exp[1]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2806));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I54 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[2]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502), .B(b_exp[2]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2851));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I55 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362), .B(b_exp[3]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2822));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I56 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[4]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504), .B(b_exp[4]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2844));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I57 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[4]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I58 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507), .A(a_exp[7]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I59 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506), .A(a_exp[6]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I60 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505), .A(a_exp[5]));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I61 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505), .B(b_exp[5]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2815));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I62 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[6]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506), .B(b_exp[6]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2838));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I63 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[7]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507), .B(b_exp[7]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2809));
INVX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I64 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10347));
INVX2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I65 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I66 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509), .A(b_exp[0]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I67 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N501), .B(b_exp[1]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2817));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I68 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N502), .B(b_exp[2]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2811));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I69 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339), .A(b_exp[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10362), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10327));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I70 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513), .A(b_exp[4]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N504), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2804));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I71 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3328), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N513), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I72 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I73 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I74 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10367));
AO22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I75 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10339), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10324), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I76 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N505), .B(b_exp[5]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2827));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I77 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N506), .B(b_exp[6]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10290));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I78 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[6]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I79 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N515), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3345));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I80 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[5]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I81 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N514), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3337));
ADDFHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I82 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N507), .B(b_exp[7]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10297));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I83 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[7]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I84 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N516), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3353));
NOR3X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I85 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10141), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10128), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10152));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I86 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[2]));
AO22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I87 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10377), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10374), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I88 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[1]));
AOI22X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I89 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[1]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3341), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N510), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]));
INVX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I90 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[1]));
INVX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I91 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
INVX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I92 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
CLKINVX12 DFT_compute_cynw_cm_float_add2_E8_M23_2_I93 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I94 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20]), .A(b_man[19]), .B(a_man[19]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MXI2XL mx2a_A_I3365 (.Y(N6856), .A(b_man[18]), .B(a_man[18]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
INVXL mx2a_A_I3366 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19]), .A(N6856));
XOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I96 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[0]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N500), .B(b_exp[0]));
AOI22X4 DFT_compute_cynw_cm_float_add2_E8_M23_2_I97 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[0]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N509), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[8]), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[0]), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3350));
CLKINVX6 DFT_compute_cynw_cm_float_add2_E8_M23_2_I98 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[0]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I99 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
MXI2XL mx2a_A_I3367 (.Y(N6863), .A(b_man[17]), .B(a_man[17]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
INVXL mx2a_A_I3368 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18]), .A(N6863));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I101 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17]), .A(b_man[16]), .B(a_man[16]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I102 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I103 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I104 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23]), .A(b_man[22]), .B(a_man[22]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I105 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I106 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22]), .A(b_man[21]), .B(a_man[21]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I107 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21]), .A(b_man[20]), .B(a_man[20]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I108 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I109 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
INVX2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I110 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I111 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
NAND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I112 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I113 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10423));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I114 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N539));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I115 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591), .A(a_man[16]), .B(b_man[16]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I116 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N591), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I117 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I118 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I119 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I120 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[19]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[18]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I121 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16]), .A(b_man[15]), .B(a_man[15]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I122 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[17]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I123 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I124 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[23]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[22]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I125 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[21]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[20]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I126 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I127 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I128 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I129 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I130 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590), .A(a_man[15]), .B(b_man[15]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I131 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N590), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I132 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3393), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I133 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I134 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15]), .A(b_man[14]), .B(a_man[14]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I135 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[16]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I136 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3503), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I137 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3481), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3414), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I138 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I139 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I140 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3535));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I141 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589), .A(a_man[14]), .B(b_man[14]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I142 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N589), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I143 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3517), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I144 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I145 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14]), .A(b_man[13]), .B(a_man[13]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I146 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[15]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I147 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I148 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3467), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I149 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3447), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3380), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I150 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I151 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I152 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3498));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I153 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588), .A(a_man[13]), .B(b_man[13]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I154 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N588), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I155 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3392));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I156 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13]), .A(b_man[12]), .B(a_man[12]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I157 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I158 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3434), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I159 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3412), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I160 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I161 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3462));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I162 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587), .A(a_man[12]), .B(b_man[12]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I163 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N587), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I164 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3516), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3534), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I165 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12]), .A(b_man[11]), .B(a_man[11]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I166 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[13]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I167 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3399), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I168 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3378), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I169 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I170 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3429));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I171 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586), .A(a_man[11]), .B(b_man[11]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I172 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N586), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I173 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3480), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3461), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I174 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11]), .A(b_man[10]), .B(a_man[10]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I175 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[12]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I176 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3525), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I177 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3502), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I178 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I179 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3394));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I180 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585), .A(a_man[10]), .B(b_man[10]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I181 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N585), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I182 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3446), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3428), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
MXI2XL mx2a_A_I3369 (.Y(N6870), .A(b_man[9]), .B(a_man[9]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
INVXL mx2a_A_I3370 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10]), .A(N6870));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3163 (.Y(N6355), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[11]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3164 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420), .A(N6355));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3165 (.Y(N6364), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3489), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3166 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487), .A(N6364));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I186 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3466), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I187 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I188 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3518));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I189 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584), .A(a_man[9]), .B(b_man[9]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I190 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N584), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I191 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9]), .A(b_man[8]), .B(a_man[8]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I192 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[10]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I193 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3454), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I194 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3433), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I195 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I196 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3482));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I197 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583), .A(a_man[8]), .B(b_man[8]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I198 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N583), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I199 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8]), .A(b_man[7]), .B(a_man[7]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I200 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[9]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I201 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3420), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I202 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3398), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I203 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3410), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I204 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3422), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I205 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[8]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3448), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I206 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[8]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I207 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582), .A(a_man[7]), .B(b_man[7]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I208 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N582), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I209 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7]), .A(b_man[6]), .B(a_man[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I210 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[8]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I211 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3387), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I212 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3523), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I213 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3376), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3418), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I214 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3476), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I215 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[7]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3413), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I216 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[7]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I217 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581), .A(a_man[6]), .B(b_man[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I218 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N581), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I219 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6]), .A(b_man[5]), .B(a_man[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I220 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I221 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3509), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I222 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3487), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I223 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3501), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3385), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I224 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3533), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I225 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[6]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3379), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I226 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[6]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I227 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580), .A(a_man[5]), .B(b_man[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I228 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N580), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I229 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5]), .A(b_man[4]), .B(a_man[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I230 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[6]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I231 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3475), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I232 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3453), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I233 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3465), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3507), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I234 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3426), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I235 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[5]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3504), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I236 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[5]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I237 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579), .A(a_man[4]), .B(b_man[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I238 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N579), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I239 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4]), .A(b_man[3]), .B(a_man[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I240 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[5]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I241 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3441), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I242 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3419), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I243 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3432), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3472), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I244 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3391), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I245 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[4]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3468), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I246 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[4]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I247 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578), .A(a_man[3]), .B(b_man[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I248 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N578), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I249 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3]), .A(b_man[2]), .B(a_man[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I250 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[4]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I251 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3406), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I252 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3405), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3386), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I253 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3397), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3438), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I254 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3515), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I255 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[3]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3435), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I256 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[3]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I257 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577), .A(a_man[2]), .B(b_man[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I258 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N577), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3167 (.Y(N6370), .A(b_man[1]), .B(a_man[1]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I3168 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2]), .A(N6370));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I260 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I261 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3531), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10346));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I262 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10363), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3508), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I263 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10369), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3521), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I264 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3479), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I265 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[2]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3400), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I266 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[2]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I267 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576), .A(a_man[1]), .B(b_man[1]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I268 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N576), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I269 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
AOI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I270 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3445), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I271 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1]), .A(b_man[0]), .B(a_man[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I272 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I273 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3496), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3425), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I274 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3495), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3474));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I275 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3485));
AOI211XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I276 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10162), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10167), .C0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10157));
NOR3X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I277 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10133), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10124), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10144));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I278 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575), .A(a_man[0]), .B(b_man[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I279 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N575), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I280 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I281 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[1]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3455));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I282 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3526), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3459), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3513), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3490));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I283 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3437), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3458), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3440), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3470));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I284 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3415), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3452), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3494), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3381));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I285 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[0]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3484), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3488), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3408), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520));
AND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I286 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N522), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[0]));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I287 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[0]));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I288 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4035));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I289 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4015));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I290 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3930));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I291 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3996));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I292 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3911));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I293 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3977));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I294 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4043));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I295 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3957));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I296 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4023));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I297 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3938));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I298 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4004));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I299 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3919));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I300 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3985));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I301 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3900));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I302 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3966));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I303 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4032));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I304 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3947));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I305 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4230), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N462));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I306 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3450));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I307 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3383));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I308 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597), .A(a_man[22]), .B(b_man[22]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I309 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N597), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I310 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3471));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I311 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596), .A(a_man[21]), .B(b_man[21]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I312 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N596), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I313 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3402));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I314 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595), .A(a_man[20]), .B(b_man[20]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I315 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N595), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I316 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3492));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I317 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594), .A(a_man[19]), .B(b_man[19]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I318 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N594), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I319 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3423));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I320 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593), .A(a_man[18]), .B(b_man[18]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I321 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N593), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
NOR4BBX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I322 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3704), .BN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3772), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3520), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3511));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I323 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592), .A(a_man[17]), .B(b_man[17]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
XNOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I324 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N592), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I325 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N420), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[1]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[1]));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I326 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N421), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[2]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4002));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I327 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N422), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[3]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3917));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I328 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N423), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[4]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[4]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3983));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I329 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N424), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[5]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[5]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4049));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I330 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N425), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[6]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[6]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3963));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I331 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N426), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[7]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4029));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I332 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N427), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[8]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[8]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3944));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I333 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N428), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[9]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[9]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4009));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I334 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N429), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[10]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[10]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3924));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I335 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N430), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[11]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[11]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3990));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I336 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N431), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[12]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[12]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3905));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I337 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N432), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[13]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[13]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3971));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I338 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N433), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[14]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4037));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I339 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N434), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[15]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[15]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3951));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I340 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N435), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[16]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[16]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4017));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I341 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N436), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[17]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[17]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3932));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I342 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N437), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3999));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I343 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N438), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3913));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I344 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N439), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3980));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I345 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N440), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4046));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I346 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N441), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3959));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I347 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N442), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4026));
ADDFX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I348 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N443), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3941));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I349 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N444));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I350 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25]));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I351 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6144), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I352 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[25]));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I353 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I354 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6150), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6149));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I355 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17]), .A0(N6124), .A1(N6007), .B0(N6073), .B1(N6122));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I356 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4206), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N461));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I357 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]), .A0(N6077), .A1(N6007), .B0(N6073), .B1(N6075));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I358 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I359 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4267), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N459));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I360 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6143), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I361 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165), .A0(N6298), .A1(N6083), .B0(N6073), .B1(N6304));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I362 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6165));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I363 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4184), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N460));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I364 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6145), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I365 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485), .A0(N6217), .A1(N6073), .B0(N6221), .B1(N6129));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I366 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N485));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I367 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I368 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I369 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4197), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N456));
INVXL buf1_A_I3391 (.Y(N6918), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4226));
INVXL buf1_A_I3392 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6152), .A(N6918));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I371 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]), .A0(N6101), .A1(N6083), .B0(N6097), .B1(N5984));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I372 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4280), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N455));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I373 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6146), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I374 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]), .A0(N6147), .A1(N6107), .B0(N6143), .B1(N5984));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I375 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I376 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4242), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N458));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I377 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483), .A0(N5984), .A1(N6228), .B0(N6230), .B1(N6129));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I378 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N483));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I379 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4220), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N457));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I380 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482), .A0(N5984), .A1(N6192), .B0(N6194), .B1(N6129));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I381 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N482));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I382 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I383 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I384 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I385 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148), .A(N6654));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I386 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25]), .A(N6185), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148));
ADDFHXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I387 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[18]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[18]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4012));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I388 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[19]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[19]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3927));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I389 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[20]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[20]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3993));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I390 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[21]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[21]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3908));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I391 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[22]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[22]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3974));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I392 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[23]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[23]), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4040));
XOR3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I393 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N469), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__39[24]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N3954));
MXI2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I394 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180), .A(N6675), .B(N6185), .S0(N6677));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3156 (.Y(N6331), .A0(N6007), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4180), .B0(N6009), .B1(N6073));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3157 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]), .A(N6331));
NOR2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I396 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I397 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4263), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N468));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I398 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493), .A0(N6253), .A1(N6073), .B0(N6257), .B1(N6007));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I399 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N493));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I400 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4239), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N467));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I401 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173), .A0(N6289), .A1(N6083), .B0(N6073), .B1(N6295));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I402 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6173));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I403 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]));
NAND2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I404 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I405 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4216), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N466));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I406 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21]), .A0(N6158), .A1(N6083), .B0(N6073), .B1(N6156));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I407 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4193), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N465));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I408 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]), .A0(N6135), .A1(N6129), .B0(N5984), .B1(N6133));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I409 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I410 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4276), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N464));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I411 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19]), .A0(N6175), .A1(N6007), .B0(N6073), .B1(N6173));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I412 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4252), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N463));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I413 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488), .A0(N5984), .A1(N6210), .B0(N6212), .B1(N6129));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I414 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N488));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I415 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I416 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338));
NOR2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I417 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411));
NAND2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I418 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I419 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4256), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N454));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I420 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479), .A0(N6073), .A1(N6262), .B0(N6266), .B1(N6107));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I421 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N479));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I422 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4234), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N453));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I423 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478), .A0(N6280), .A1(N6073), .B0(N6284), .B1(N6107));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I424 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N478));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I425 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I426 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4210), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N452));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I427 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477), .A0(N6271), .A1(N6073), .B0(N6275), .B1(N6107));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I428 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N477));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I429 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4188), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N451));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3159 (.Y(N6341), .A0(N6113), .A1(N6107), .B0(N6109), .B1(N5984));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3160 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]), .A(N6341));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I431 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I432 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I433 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4271), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N450));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I434 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6147), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6142));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I435 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475), .A0(N5984), .A1(N6246), .B0(N6248), .B1(N5981));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I436 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N475));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I437 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4247), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N449));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I438 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474), .A0(N5984), .A1(N6201), .B0(N6203), .B1(N5981));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I439 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N474));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I440 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I441 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4224), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N448));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I442 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473), .A0(N6235), .A1(N5984), .B0(N6239), .B1(N5981));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I443 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N473));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I444 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4200), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N447));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3161 (.Y(N6349), .A0(N6089), .A1(N6083), .B0(N5984), .B1(N6087));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I3162 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]), .A(N6349));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I446 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I447 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I448 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I449 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4380), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I450 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I451 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4411), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4354), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4374));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I452 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4420), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4393));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I453 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I454 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I455 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6212));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I456 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4412), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4336));
OAI2BB1X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I457 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376), .A0N(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4345), .A1N(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4384), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4364));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I458 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4375), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4395));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I459 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4426));
AOI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I460 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4405), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4415), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4339));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I461 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4338), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4359));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I462 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4388));
AOI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I463 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4366), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4348), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4367));
AOI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I464 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4360), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4389));
OA21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I465 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4376), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4342));
BUFX3 DFT_compute_cynw_cm_float_add2_E8_M23_2_I466 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I467 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I468 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I469 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21]));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I470 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4370), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4392));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I471 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I472 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25]));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I473 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4400), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4423));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I474 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4335), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4414), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4347));
INVX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I475 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I476 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I477 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I478 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4408), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4428));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I479 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I480 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17]));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I481 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4341), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4362));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I482 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4355), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4401), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4383));
NAND2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I483 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372));
NAND2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I484 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10223), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10211));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I485 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4259), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N445));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I486 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470), .A0(N5984), .A1(N5977), .B0(N5979), .B1(N5981));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I487 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N470));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I488 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4177), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[24]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__55[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N446));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I489 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471), .A0(N5984), .A1(N5986), .B0(N5988), .B1(N5981));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I490 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N471));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I491 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]));
NOR2X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I492 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4352));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I493 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I494 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I495 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4349), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4368));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I496 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I497 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]));
OAI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I498 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4378), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4398));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I499 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4371), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4390), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4421));
AOI21X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I500 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10217), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10220));
NOR2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I501 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417));
NOR2X2 DFT_compute_cynw_cm_float_add2_E8_M23_2_I502 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10221), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10208));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I503 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I504 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4775));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I505 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I506 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I507 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I508 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4402), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4407));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I509 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372));
AOI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I510 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4418), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4382), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4404));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I511 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3]));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I512 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I513 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[22]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I514 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I515 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4779), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I516 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I517 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[21]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I518 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4741), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I519 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I520 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I521 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I522 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[24]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I523 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4852), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I524 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I525 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[23]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I526 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4818), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I527 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4803), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I528 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4742), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I529 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I530 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[18]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I531 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4799), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I532 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I533 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[17]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I534 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4763), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I535 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I536 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I537 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[20]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I538 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4875), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I539 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I540 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[19]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I541 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4836), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I542 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I543 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I544 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I545 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[24]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4796), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I546 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N498), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I547 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I548 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I549 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I550 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
AND4XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I551 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[4]), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I552 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I553 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4593), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4603), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[6]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I554 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I555 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
NAND3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I556 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205), .A(N4572), .B(N5467), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[25]));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I557 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499), .A(N5139), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6205));
OR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I558 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .A(N4892), .B(N4894), .C(N3881), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N499));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I559 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4351));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I560 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[3]));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I561 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570), .A(N5154), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I562 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573), .A(N5467), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I563 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[0]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10019), .B(b_exp[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2914));
AOI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I564 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10197), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4372), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10202));
OAI21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I565 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[0]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4417), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10209), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10216));
NAND2BXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I566 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578), .AN(N5508), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[0]));
OAI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I567 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4573), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4578), .B0(N5467), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I568 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4571), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]));
OR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I569 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557), .A(N5409), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2]));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I570 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4561), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4557), .B0(N5409), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[2]));
OAI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I571 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4570), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4567), .B0(N5154), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I572 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566), .A(N6657));
OR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I573 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]));
AOI22X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I574 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4575), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4554), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4566), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]));
NOR4X1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I575 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73), .A(N4038), .B(N6666), .C(N4572), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4552));
NOR4X6 DFT_compute_cynw_cm_float_add2_E8_M23_2_I576 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72), .A(N4293), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5]), .D(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__73));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I577 (.Y(x[22]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[24]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I578 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4863), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4825), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I579 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4766), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4728), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I580 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4876), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I581 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[0]));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I582 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[8]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[16]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I583 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[4]), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4895), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I584 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4884), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I585 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4787), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4749), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I586 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I587 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[23]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4759), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I588 (.Y(x[21]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[23]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I589 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4765), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4837), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I590 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[7]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[15]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I591 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4859), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I592 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4846), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I593 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4861), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I594 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[22]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4893), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I595 (.Y(x[20]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[22]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I596 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4898), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4801), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I597 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[6]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[14]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I598 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4822), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I599 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4772), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I600 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4823), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I601 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[21]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4855), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I602 (.Y(x[19]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[21]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I603 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[5]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[13]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I604 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4784), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I605 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4870), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I606 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4786), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I607 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[20]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4820), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I608 (.Y(x[18]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[20]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I609 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[4]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[12]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I610 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4746), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I611 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4794), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I612 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4748), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I613 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[19]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4781), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I614 (.Y(x[17]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[19]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I615 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[11]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I616 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4881), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I617 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4890), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I618 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4883), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I619 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[18]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4744), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I620 (.Y(x[16]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[18]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I621 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[10]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I622 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4842), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I623 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4817), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I624 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4845), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I625 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[17]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4878), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I626 (.Y(x[15]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[17]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I627 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[1]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__51[9]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4867));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I628 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4807), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I629 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4740), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I630 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4809), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I631 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[16]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4840), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I632 (.Y(x[14]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[16]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I633 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4769), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I634 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4835), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I635 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4770), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I636 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[15]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4804), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I637 (.Y(x[13]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[15]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I638 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4866), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I639 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4762), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I640 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4733), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I641 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[14]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4767), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I642 (.Y(x[12]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[14]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I643 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4790), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I644 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4858), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I645 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4869), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I646 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[13]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4729), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I647 (.Y(x[11]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[13]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I648 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4887), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I649 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4783), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I650 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4830), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I651 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[12]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4864), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I652 (.Y(x[10]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[12]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I653 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4814), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I654 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4880), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I655 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4793), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I656 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[11]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4826), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I657 (.Y(x[9]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[11]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I658 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4736), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I659 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4806), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I660 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4753), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I661 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[10]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4788), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I662 (.Y(x[8]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[10]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I663 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4833), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I664 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4731), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I665 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4888), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I666 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[9]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4750), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I667 (.Y(x[7]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[9]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I668 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4760), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I669 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4828), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I670 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4851), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I671 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[8]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4885), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I672 (.Y(x[6]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[8]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I673 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4856), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I674 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4752), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4897));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I675 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4816), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I676 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[7]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4847), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I677 (.Y(x[5]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[7]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I678 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4844), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4849));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I679 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4812), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4778), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I680 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[6]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4811), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I681 (.Y(x[4]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I682 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4739), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I683 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[5]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4773), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4755), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I684 (.Y(x[3]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NAND2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I685 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4798), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6154));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I686 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[4]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6161), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4734), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4853), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I687 (.Y(x[2]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I688 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[3]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4871));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I689 (.Y(x[1]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
NOR2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I690 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[2]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4758), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4831));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I691 (.Y(x[0]), .A(N6854), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I692 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I693 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654), .A(N6666));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I694 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4644), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[2]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1]));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I695 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4632), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4668), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[3]), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4657));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I696 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639), .A(N6657), .B(N6663));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I697 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4660), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[5]));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I698 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4652), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__40[1]));
ADDHX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I699 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[0]), .A(N5508), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4645));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I700 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[1]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4569), .B(N5475), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4653));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I701 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[2]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4640), .B(N5398), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4646));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I702 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[3]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4565), .B(N5145), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4670));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I703 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[4]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4635), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4639), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4641));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I704 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[5]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4650), .B(N4578), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4662));
ADDFXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I705 (.CO(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655), .S(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[6]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4654), .B(N4572), .CI(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4636));
XNOR3XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I706 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[7]), .A(N4038), .B(N6666), .C(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4655));
AO22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I707 (.Y(x[30]), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6216), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[7]), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I708 (.Y(x[29]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[6]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I709 (.Y(x[28]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[5]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I710 (.Y(x[27]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[4]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I711 (.Y(x[26]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[3]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I712 (.Y(x[25]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[2]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I713 (.Y(x[24]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[1]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
MX2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I714 (.Y(x[23]), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__77), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__66[0]), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__72));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I715 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10111));
INVXL DFT_compute_cynw_cm_float_add2_E8_M23_2_I716 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888), .A(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N10417));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I717 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4159), .A0(b_sign), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888), .B0(a_sign), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I718 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418), .AN(a_sign), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__28));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I719 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417), .AN(b_sign), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__31));
AOI22XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I720 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N4164), .A0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N418), .A1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2888), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N417), .B1(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N2842));
MXI2XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I721 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52), .A(N4903), .B(N4901), .S0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N6148));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I722 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__52), .B(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[5]));
AO21XL DFT_compute_cynw_cm_float_add2_E8_M23_2_I723 (.Y(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69), .A0(N4247), .A1(N4249), .B0(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_N496));
NOR2BX1 DFT_compute_cynw_cm_float_add2_E8_M23_2_I724 (.Y(x[31]), .AN(DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__69), .B(N6854));
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__44[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[2] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[4] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[5] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[6] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__47[7] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__48[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[9] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[10] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[11] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[12] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[13] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[14] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[15] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[16] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[17] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[18] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[19] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[20] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[21] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[22] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[23] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__49[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_delta[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[1] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[2] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[3] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[4] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[5] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[6] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[7] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[8] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[9] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[10] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[11] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[12] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[13] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[14] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[15] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[16] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[17] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[18] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[19] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[20] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[21] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[22] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[23] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__56[24] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[0] = 1'B0;
assign DFT_compute_cynw_cm_float_add2_E8_M23_1_inst_inst_cellmath__63[1] = 1'B0;
endmodule

/* CADENCE  ubn4SA7dohw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



