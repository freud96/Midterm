/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:22:23 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_mul_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire  inst_cellmath__17,
	inst_cellmath__18,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23,
	inst_cellmath__24,
	inst_cellmath__25,
	inst_cellmath__26,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__32,
	inst_cellmath__33;
wire [9:0] inst_cellmath__34;
wire  inst_cellmath__37,
	inst_cellmath__38,
	inst_cellmath__41,
	inst_cellmath__42;
wire [47:0] inst_cellmath__43;
wire [7:0] inst_cellmath__50,
	inst_cellmath__54;
wire  inst_cellmath__56,
	inst_cellmath__60,
	inst_cellmath__61;
wire N267,N268,N269,N270,N272,N273,N274 
	,N276,N1314,N1318,N1338,N1340,N1361,N1369,N1372 
	,N1374,N1378,N1380,N1383,N1389,N1393,N1425,N1429 
	,N1449,N1451,N1472,N1480,N1483,N1485,N1489,N1491 
	,N1494,N1500,N1504,N1551,N1552,N1553,N1554,N1555 
	,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563 
	,N1564,N1566,N1567,N1568,N1569,N1570,N1571,N1572 
	,N1574,N1576,N1577,N1578,N1579,N1580,N1581,N1582 
	,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590 
	,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1599 
	,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607 
	,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1616 
	,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624 
	,N1625,N1626,N1627,N1628,N1630,N1631,N1632,N1633 
	,N1634,N1636,N1637,N1638,N1639,N1640,N1641,N1642 
	,N1643,N1644,N1645,N1646,N1647,N1648,N1650,N1651 
	,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659 
	,N1660,N1661,N1662,N1664,N1665,N1666,N1667,N1668 
	,N1669,N1670,N1671,N1673,N1674,N1675,N1676,N1677 
	,N1678,N1679,N1680,N1681,N1683,N1684,N1685,N1686 
	,N1687,N1689,N1690,N1691,N1692,N1693,N1694,N1695 
	,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703 
	,N1704,N1705,N1707,N1708,N1709,N1710,N1711,N1712 
	,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720 
	,N1721,N1722,N1723,N1725,N1726,N1727,N1728,N1729 
	,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737 
	,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745 
	,N1746,N1747,N1748,N1750,N1751,N1752,N1753,N1754 
	,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762 
	,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1771 
	,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780 
	,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788 
	,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798 
	,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806 
	,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814 
	,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822 
	,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1832 
	,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840 
	,N1841,N1842,N1843,N1844,N1845,N1847,N1848,N1849 
	,N1851,N1852,N1853,N1854,N1855,N1856,N1858,N1859 
	,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867 
	,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875 
	,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883 
	,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891 
	,N1892,N1893,N1894,N1896,N1897,N1898,N1899,N1900 
	,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908 
	,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916 
	,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925 
	,N1926,N1927,N1929,N1930,N1931,N1932,N1933,N1934 
	,N1935,N1936,N1938,N1939,N1940,N1942,N1943,N1944 
	,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952 
	,N1953,N1954,N1956,N1957,N1958,N1959,N1960,N1961 
	,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969 
	,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978 
	,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986 
	,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994 
	,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2003 
	,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011 
	,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019 
	,N2020,N2022,N2023,N2024,N2025,N2026,N2027,N2028 
	,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036 
	,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044 
	,N2045,N2046,N2047,N2048,N2049,N2051,N2052,N2053 
	,N2054,N2055,N2056,N2057,N2058,N2060,N2061,N2062 
	,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071 
	,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080 
	,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2089 
	,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097 
	,N2098,N2100,N2101,N2102,N2103,N2104,N2105,N2106 
	,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115 
	,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123 
	,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131 
	,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139 
	,N2140,N2141,N2142,N2143,N2144,N2145,N2147,N2148 
	,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156 
	,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164 
	,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172 
	,N2173,N2174,N2175,N2176,N2177,N2179,N2180,N2181 
	,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189 
	,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197 
	,N2198,N2199,N2200,N2203,N2204,N2205,N2206,N2207 
	,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215 
	,N2216,N2217,N2219,N2220,N2221,N2222,N2223,N2224 
	,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2233 
	,N2234,N2235,N2236,N2238,N2239,N2240,N2241,N2242 
	,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250 
	,N2251,N2253,N2254,N2255,N2256,N2257,N2258,N2259 
	,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267 
	,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2276 
	,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284 
	,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292 
	,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300 
	,N2301,N2302,N2303,N2304,N2305,N2306,N2308,N2309 
	,N2310,N2311,N2313,N2314,N2315,N2317,N2318,N2319 
	,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2328 
	,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336 
	,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344 
	,N2345,N2346,N2347,N2348,N2350,N2352,N2353,N2355 
	,N2356,N2357,N2358,N2360,N2361,N2362,N2363,N2364 
	,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372 
	,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380 
	,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389 
	,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397 
	,N2398,N2400,N2401,N2402,N2403,N2404,N2405,N2406 
	,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414 
	,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422 
	,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430 
	,N2431,N2432,N2434,N2435,N2436,N2437,N2438,N2439 
	,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447 
	,N2448,N2449,N2450,N2451,N2452,N2454,N2455,N2456 
	,N2457,N2459,N2460,N2461,N2463,N2464,N2465,N2466 
	,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474 
	,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482 
	,N2483,N2484,N2485,N2486,N2487,N2488,N2490,N2491 
	,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499 
	,N2500,N2501,N2502,N2503,N2505,N2506,N2507,N2508 
	,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516 
	,N2517,N2518,N2519,N2521,N2522,N2523,N2524,N2525 
	,N2526,N2527,N2529,N2531,N2532,N2533,N2534,N2535 
	,N2536,N2537,N2538,N2540,N2541,N2542,N2543,N2544 
	,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552 
	,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560 
	,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568 
	,N2569,N2570,N2571,N2572,N2574,N2575,N2576,N2577 
	,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586 
	,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594 
	,N2595,N2596,N2597,N2598,N2600,N2601,N2602,N2603 
	,N2604,N2605,N2606,N2608,N2610,N2611,N2612,N2613 
	,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621 
	,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629 
	,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638 
	,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646 
	,N2647,N2648,N2650,N2651,N2652,N2653,N2654,N2655 
	,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663 
	,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671 
	,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679 
	,N2680,N2681,N2683,N2684,N2685,N2686,N2687,N2688 
	,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696 
	,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704 
	,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714 
	,N2715,N2716,N2717,N2719,N2721,N2722,N2723,N2724 
	,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732 
	,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740 
	,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748 
	,N2749,N2750,N2751,N2752,N2754,N2755,N2756,N2757 
	,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765 
	,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773 
	,N2774,N2775,N2776,N2778,N2779,N2780,N2781,N2782 
	,N2783,N2784,N2785,N2786,N2788,N2789,N2790,N2791 
	,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799 
	,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807 
	,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815 
	,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823 
	,N2824,N2825,N2827,N2828,N2829,N2830,N2832,N2833 
	,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841 
	,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849 
	,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857 
	,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2867 
	,N2868,N2869,N2871,N2872,N2873,N2874,N2875,N2876 
	,N2877,N2878,N2879,N2880,N2882,N2883,N2884,N2885 
	,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893 
	,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901 
	,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909 
	,N2910,N2911,N2913,N2914,N2915,N2916,N2917,N2918 
	,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926 
	,N2927,N2928,N2930,N2931,N2932,N2933,N2934,N2935 
	,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2944 
	,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952 
	,N2953,N2955,N2956,N2957,N2958,N2959,N2961,N2962 
	,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970 
	,N2971,N2972,N2973,N2974,N2975,N2976,N2978,N2979 
	,N2980,N2981,N2982,N2983,N2985,N2986,N2987,N2988 
	,N2989,N2990,N2991,N2993,N2994,N2995,N2996,N2997 
	,N2998,N2999,N3000,N3001,N3003,N3004,N3005,N3006 
	,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014 
	,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022 
	,N3023,N3025,N3026,N3027,N3028,N3029,N3030,N3031 
	,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040 
	,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048 
	,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3057 
	,N3058,N3059,N3061,N3062,N3063,N3064,N3065,N3066 
	,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3075 
	,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083 
	,N3084,N3086,N3087,N3088,N3089,N3090,N3091,N3092 
	,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100 
	,N3101,N3102,N3103,N3104,N3105,N3107,N3108,N3109 
	,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117 
	,N3118,N3119,N3120,N3121,N3122,N3124,N3125,N3126 
	,N3127,N3128,N3130,N3131,N3133,N3134,N3135,N3136 
	,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144 
	,N3145,N3146,N3147,N3149,N3150,N3151,N3152,N3153 
	,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161 
	,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169 
	,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177 
	,N3178,N3179,N3181,N3182,N3183,N3184,N3185,N3186 
	,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194 
	,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3203 
	,N3205,N3206,N3208,N3209,N3210,N3211,N3212,N3213 
	,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222 
	,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230 
	,N3231,N3232,N3233,N3234,N3235,N3237,N3238,N3239 
	,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247 
	,N3248,N3249,N3250,N3251,N3252,N3253,N3255,N3256 
	,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264 
	,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272 
	,N3273,N3274,N3275,N3276,N3277,N3279,N3280,N3281 
	,N3282,N3283,N3284,N3285,N3286,N3288,N3289,N3290 
	,N3291,N3292,N3293,N3295,N3296,N3297,N3298,N3299 
	,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307 
	,N3308,N3309,N3310,N3312,N3313,N3314,N3315,N3316 
	,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324 
	,N3325,N3327,N3328,N3329,N3330,N3331,N3332,N3333 
	,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341 
	,N3342,N3343,N3344,N3345,N3346,N3348,N3349,N3350 
	,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358 
	,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367 
	,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375 
	,N3376,N3377,N3378,N3379,N3380,N3381,N3384,N3385 
	,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3395 
	,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403 
	,N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411 
	,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419 
	,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427 
	,N3428,N3429,N3430,N3431,N3433,N3434,N3435,N3436 
	,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444 
	,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453 
	,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461 
	,N3462,N3464,N3465,N3466,N3467,N3468,N3469,N3470 
	,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478 
	,N3479,N3480,N3481,N3482,N3483,N3485,N3486,N3487 
	,N3488,N3489,N3490,N3491,N3492,N3493,N3495,N3496 
	,N3497,N3498,N3499,N3500,N3501,N3502,N3504,N3505 
	,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N5430 
	,N5437,N5449,N5452,N5456,N5457,N5462,N5468,N5472 
	,N5477,N5480,N5501,N5505,N5507,N5529,N5530,N5534 
	,N5538,N5564,N5566,N5575,N5580,N5618,N5620,N5622 
	,N5625,N5627,N5631,N5633,N5641,N5669,N5672,N5673 
	,N5677,N5680,N5682,N5684,N5687,N5692,N5694,N5697 
	,N5700,N5701,N5705,N5707,N5711,N5714,N5719,N5722 
	,N5727,N5729,N5732,N5735,N5741,N5743,N5747,N5750 
	,N5755,N5759,N5762,N5766,N5767,N5770,N5776,N5778 
	,N8064,N8072,N8078,N8085,N16704;
XOR2XL cynw_cm_float_mul_I195 (.Y(inst_cellmath__33), .A(a_sign), .B(b_sign));
OR4X1 inst_cellmath__26__8__I9644 (.Y(N1314), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__26__8__I9645 (.Y(N1318), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL inst_cellmath__26__8__I202 (.Y(inst_cellmath__26), .A(N1314), .B(N1318));
NAND2XL inst_cellmath__17_0_I203 (.Y(N1338), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__17_0_I9646 (.Y(N1340), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3440 (.Y(N8064), .A(a_exp[7]), .B(a_exp[6]), .C(N1340));
NOR2XL hyperpropagate_4_1_A_I3441 (.Y(inst_cellmath__17), .A(N1338), .B(N8064));
NOR2XL inst_cellmath__19__5__I216 (.Y(N1361), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__19__5__I217 (.Y(N1369), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__19__5__I218 (.Y(N1380), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__19__5__I219 (.Y(N1389), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__19__5__I9647 (.Y(N1374), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__19__5__I9648 (.Y(N1383), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__19__5__I9649 (.Y(N1393), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__19__5__I223 (.Y(N1378), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N1374));
NAND4XL inst_cellmath__19__5__I225 (.Y(N1372), .A(N1361), .B(N1380), .C(N1369), .D(N1389));
NOR4BX1 inst_cellmath__19__5__I9650 (.Y(inst_cellmath__19), .AN(N1378), .B(N1372), .C(N1383), .D(N1393));
AND2XL cynw_cm_float_mul_I228 (.Y(inst_cellmath__23), .A(inst_cellmath__17), .B(inst_cellmath__19));
AND2XL cynw_cm_float_mul_I229 (.Y(N268), .A(inst_cellmath__26), .B(inst_cellmath__23));
OR4X1 inst_cellmath__25__7__I9651 (.Y(N1425), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__25__7__I9652 (.Y(N1429), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__25__7__I236 (.Y(inst_cellmath__25), .A(N1425), .B(N1429));
NAND2XL inst_cellmath__18_0_I237 (.Y(N1449), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__18_0_I9653 (.Y(N1451), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3442 (.Y(N8072), .A(b_exp[7]), .B(b_exp[6]), .C(N1451));
NOR2XL hyperpropagate_4_1_A_I3443 (.Y(inst_cellmath__18), .A(N1449), .B(N8072));
NOR2XL inst_cellmath__20__6__I250 (.Y(N1472), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__20__6__I251 (.Y(N1480), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__20__6__I252 (.Y(N1491), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__20__6__I253 (.Y(N1500), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__20__6__I9654 (.Y(N1485), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__20__6__I9655 (.Y(N1494), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__20__6__I9656 (.Y(N1504), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__20__6__I257 (.Y(N1489), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N1485));
NAND4XL inst_cellmath__20__6__I259 (.Y(N1483), .A(N1472), .B(N1491), .C(N1480), .D(N1500));
NOR4BX1 inst_cellmath__20__6__I9657 (.Y(inst_cellmath__20), .AN(N1489), .B(N1483), .C(N1494), .D(N1504));
AND2XL cynw_cm_float_mul_I262 (.Y(inst_cellmath__24), .A(inst_cellmath__18), .B(inst_cellmath__20));
AND2XL cynw_cm_float_mul_I263 (.Y(N267), .A(inst_cellmath__25), .B(inst_cellmath__24));
NOR2BX1 cynw_cm_float_mul_I264 (.Y(inst_cellmath__21), .AN(inst_cellmath__17), .B(inst_cellmath__19));
NOR2BX1 cynw_cm_float_mul_I265 (.Y(inst_cellmath__22), .AN(inst_cellmath__18), .B(inst_cellmath__20));
OR4X1 cynw_cm_float_mul_I266 (.Y(inst_cellmath__29), .A(inst_cellmath__22), .B(inst_cellmath__21), .C(N268), .D(N267));
NOR2BX1 cynw_cm_float_mul_I267 (.Y(x[31]), .AN(inst_cellmath__33), .B(inst_cellmath__29));
INVXL inst_cellmath__43_0_I268 (.Y(N3303), .A(b_man[0]));
INVXL inst_cellmath__43_0_I269 (.Y(N1765), .A(b_man[1]));
INVXL inst_cellmath__43_0_I270 (.Y(N2196), .A(b_man[2]));
INVXL inst_cellmath__43_0_I271 (.Y(N2623), .A(b_man[3]));
INVXL inst_cellmath__43_0_I272 (.Y(N3050), .A(b_man[4]));
INVXL inst_cellmath__43_0_I273 (.Y(N3477), .A(b_man[5]));
INVXL inst_cellmath__43_0_I274 (.Y(N1948), .A(b_man[6]));
INVXL inst_cellmath__43_0_I275 (.Y(N2375), .A(b_man[7]));
INVXL inst_cellmath__43_0_I276 (.Y(N2806), .A(b_man[8]));
INVXL inst_cellmath__43_0_I277 (.Y(N3228), .A(b_man[9]));
INVXL inst_cellmath__43_0_I278 (.Y(N1702), .A(b_man[10]));
INVXL inst_cellmath__43_0_I279 (.Y(N2122), .A(b_man[11]));
INVXL inst_cellmath__43_0_I280 (.Y(N2556), .A(b_man[12]));
INVXL inst_cellmath__43_0_I281 (.Y(N2978), .A(b_man[13]));
INVXL inst_cellmath__43_0_I282 (.Y(N3412), .A(b_man[14]));
INVXL inst_cellmath__43_0_I283 (.Y(N1871), .A(b_man[15]));
INVXL inst_cellmath__43_0_I284 (.Y(N2301), .A(b_man[16]));
INVXL inst_cellmath__43_0_I285 (.Y(N2729), .A(b_man[17]));
INVXL inst_cellmath__43_0_I286 (.Y(N3157), .A(b_man[18]));
INVXL inst_cellmath__43_0_I287 (.Y(N1623), .A(b_man[19]));
INVXL inst_cellmath__43_0_I288 (.Y(N2049), .A(b_man[20]));
INVXL inst_cellmath__43_0_I289 (.Y(N2480), .A(b_man[21]));
INVXL inst_cellmath__43_0_I290 (.Y(N2905), .A(b_man[22]));
INVXL inst_cellmath__43_0_I291 (.Y(N3335), .A(a_man[0]));
NOR2XL inst_cellmath__43_0_I294 (.Y(N3452), .A(N3335), .B(N2196));
NOR2XL inst_cellmath__43_0_I295 (.Y(N2347), .A(N3335), .B(N2623));
NOR2XL inst_cellmath__43_0_I296 (.Y(N3201), .A(N3335), .B(N3050));
NOR2XL inst_cellmath__43_0_I297 (.Y(N2096), .A(N3335), .B(N3477));
NOR2XL inst_cellmath__43_0_I298 (.Y(N2951), .A(N3335), .B(N1948));
NOR2XL inst_cellmath__43_0_I299 (.Y(N1845), .A(N3335), .B(N2375));
NOR2XL inst_cellmath__43_0_I300 (.Y(N2701), .A(N3335), .B(N2806));
NOR2XL inst_cellmath__43_0_I301 (.Y(N1596), .A(N3335), .B(N3228));
NOR2XL inst_cellmath__43_0_I302 (.Y(N2452), .A(N3335), .B(N1702));
NOR2XL inst_cellmath__43_0_I303 (.Y(N3308), .A(N3335), .B(N2122));
NOR2XL inst_cellmath__43_0_I304 (.Y(N2199), .A(N3335), .B(N2556));
NOR2XL inst_cellmath__43_0_I305 (.Y(N3055), .A(N3335), .B(N2978));
NOR2XL inst_cellmath__43_0_I306 (.Y(N1952), .A(N3335), .B(N3412));
NOR2XL inst_cellmath__43_0_I307 (.Y(N2810), .A(N3335), .B(N1871));
NOR2XL inst_cellmath__43_0_I308 (.Y(N1705), .A(N3335), .B(N2301));
NOR2XL inst_cellmath__43_0_I309 (.Y(N2562), .A(N3335), .B(N2729));
NOR2XL inst_cellmath__43_0_I310 (.Y(N3415), .A(N3335), .B(N3157));
NOR2XL inst_cellmath__43_0_I311 (.Y(N2306), .A(N3335), .B(N1623));
NOR2XL inst_cellmath__43_0_I312 (.Y(N3164), .A(N3335), .B(N2049));
NOR2XL inst_cellmath__43_0_I313 (.Y(N2053), .A(N3335), .B(N2480));
NOR2XL inst_cellmath__43_0_I314 (.Y(N2911), .A(N3335), .B(N2905));
INVXL inst_cellmath__43_0_I315 (.Y(N1806), .A(N3335));
INVXL inst_cellmath__43_0_I316 (.Y(N1798), .A(a_man[1]));
NOR2XL inst_cellmath__43_0_I318 (.Y(N2339), .A(N1798), .B(N1765));
NOR2XL inst_cellmath__43_0_I319 (.Y(N3194), .A(N1798), .B(N2196));
NOR2XL inst_cellmath__43_0_I320 (.Y(N2086), .A(N1798), .B(N2623));
NOR2XL inst_cellmath__43_0_I321 (.Y(N2942), .A(N1798), .B(N3050));
NOR2XL inst_cellmath__43_0_I322 (.Y(N1837), .A(N1798), .B(N3477));
NOR2XL inst_cellmath__43_0_I323 (.Y(N2693), .A(N1798), .B(N1948));
NOR2XL inst_cellmath__43_0_I324 (.Y(N1588), .A(N1798), .B(N2375));
NOR2XL inst_cellmath__43_0_I325 (.Y(N2446), .A(N1798), .B(N2806));
NOR2XL inst_cellmath__43_0_I326 (.Y(N3298), .A(N1798), .B(N3228));
NOR2XL inst_cellmath__43_0_I327 (.Y(N2190), .A(N1798), .B(N1702));
NOR2XL inst_cellmath__43_0_I328 (.Y(N3044), .A(N1798), .B(N2122));
NOR2XL inst_cellmath__43_0_I329 (.Y(N1942), .A(N1798), .B(N2556));
NOR2XL inst_cellmath__43_0_I330 (.Y(N2799), .A(N1798), .B(N2978));
NOR2XL inst_cellmath__43_0_I331 (.Y(N1696), .A(N1798), .B(N3412));
NOR2XL inst_cellmath__43_0_I332 (.Y(N2551), .A(N1798), .B(N1871));
NOR2XL inst_cellmath__43_0_I333 (.Y(N3406), .A(N1798), .B(N2301));
NOR2XL inst_cellmath__43_0_I334 (.Y(N2296), .A(N1798), .B(N2729));
NOR2XL inst_cellmath__43_0_I335 (.Y(N3153), .A(N1798), .B(N3157));
NOR2XL inst_cellmath__43_0_I336 (.Y(N2041), .A(N1798), .B(N1623));
NOR2XL inst_cellmath__43_0_I337 (.Y(N2901), .A(N1798), .B(N2049));
NOR2XL inst_cellmath__43_0_I338 (.Y(N1794), .A(N1798), .B(N2480));
NOR2XL inst_cellmath__43_0_I339 (.Y(N2652), .A(N1798), .B(N2905));
INVXL inst_cellmath__43_0_I340 (.Y(N3508), .A(N1798));
INVXL inst_cellmath__43_0_I341 (.Y(N2408), .A(a_man[2]));
NOR2XL inst_cellmath__43_0_I342 (.Y(N3184), .A(N2408), .B(N3303));
NOR2XL inst_cellmath__43_0_I343 (.Y(N2077), .A(N2408), .B(N1765));
NOR2XL inst_cellmath__43_0_I344 (.Y(N2932), .A(N2408), .B(N2196));
NOR2XL inst_cellmath__43_0_I345 (.Y(N1827), .A(N2408), .B(N2623));
NOR2XL inst_cellmath__43_0_I346 (.Y(N2685), .A(N2408), .B(N3050));
NOR2XL inst_cellmath__43_0_I347 (.Y(N1578), .A(N2408), .B(N3477));
NOR2XL inst_cellmath__43_0_I348 (.Y(N2437), .A(N2408), .B(N1948));
NOR2XL inst_cellmath__43_0_I349 (.Y(N3290), .A(N2408), .B(N2375));
NOR2XL inst_cellmath__43_0_I350 (.Y(N2181), .A(N2408), .B(N2806));
NOR2XL inst_cellmath__43_0_I351 (.Y(N3035), .A(N2408), .B(N3228));
NOR2XL inst_cellmath__43_0_I352 (.Y(N1932), .A(N2408), .B(N1702));
NOR2XL inst_cellmath__43_0_I353 (.Y(N2790), .A(N2408), .B(N2122));
NOR2XL inst_cellmath__43_0_I354 (.Y(N1685), .A(N2408), .B(N2556));
NOR2XL inst_cellmath__43_0_I355 (.Y(N2543), .A(N2408), .B(N2978));
NOR2XL inst_cellmath__43_0_I356 (.Y(N3397), .A(N2408), .B(N3412));
NOR2XL inst_cellmath__43_0_I357 (.Y(N2288), .A(N2408), .B(N1871));
NOR2XL inst_cellmath__43_0_I358 (.Y(N3144), .A(N2408), .B(N2301));
NOR2XL inst_cellmath__43_0_I359 (.Y(N2032), .A(N2408), .B(N2729));
NOR2XL inst_cellmath__43_0_I360 (.Y(N2893), .A(N2408), .B(N3157));
NOR2XL inst_cellmath__43_0_I361 (.Y(N1784), .A(N2408), .B(N1623));
NOR2XL inst_cellmath__43_0_I362 (.Y(N2641), .A(N2408), .B(N2049));
NOR2XL inst_cellmath__43_0_I363 (.Y(N3498), .A(N2408), .B(N2480));
NOR2XL inst_cellmath__43_0_I364 (.Y(N2393), .A(N2408), .B(N2905));
INVXL inst_cellmath__43_0_I365 (.Y(N3247), .A(N2408));
INVXL inst_cellmath__43_0_I366 (.Y(N2835), .A(a_man[3]));
NOR2XL inst_cellmath__43_0_I367 (.Y(N2923), .A(N2835), .B(N3303));
NOR2XL inst_cellmath__43_0_I368 (.Y(N1817), .A(N2835), .B(N1765));
NOR2XL inst_cellmath__43_0_I369 (.Y(N2675), .A(N2835), .B(N2196));
NOR2XL inst_cellmath__43_0_I370 (.Y(N1567), .A(N2835), .B(N2623));
NOR2XL inst_cellmath__43_0_I371 (.Y(N2427), .A(N2835), .B(N3050));
NOR2XL inst_cellmath__43_0_I372 (.Y(N3280), .A(N2835), .B(N3477));
NOR2XL inst_cellmath__43_0_I373 (.Y(N2173), .A(N2835), .B(N1948));
NOR2XL inst_cellmath__43_0_I374 (.Y(N3027), .A(N2835), .B(N2375));
NOR2XL inst_cellmath__43_0_I375 (.Y(N1922), .A(N2835), .B(N2806));
NOR2XL inst_cellmath__43_0_I376 (.Y(N2780), .A(N2835), .B(N3228));
NOR2XL inst_cellmath__43_0_I377 (.Y(N1675), .A(N2835), .B(N1702));
NOR2XL inst_cellmath__43_0_I378 (.Y(N2534), .A(N2835), .B(N2122));
NOR2XL inst_cellmath__43_0_I379 (.Y(N3387), .A(N2835), .B(N2556));
NOR2XL inst_cellmath__43_0_I380 (.Y(N2278), .A(N2835), .B(N2978));
NOR2XL inst_cellmath__43_0_I381 (.Y(N3135), .A(N2835), .B(N3412));
NOR2XL inst_cellmath__43_0_I382 (.Y(N2024), .A(N2835), .B(N1871));
NOR2XL inst_cellmath__43_0_I383 (.Y(N2884), .A(N2835), .B(N2301));
NOR2XL inst_cellmath__43_0_I384 (.Y(N1776), .A(N2835), .B(N2729));
NOR2XL inst_cellmath__43_0_I385 (.Y(N2634), .A(N2835), .B(N3157));
NOR2XL inst_cellmath__43_0_I386 (.Y(N3486), .A(N2835), .B(N1623));
NOR2XL inst_cellmath__43_0_I387 (.Y(N2386), .A(N2835), .B(N2049));
NOR2XL inst_cellmath__43_0_I388 (.Y(N3239), .A(N2835), .B(N2480));
NOR2XL inst_cellmath__43_0_I389 (.Y(N2134), .A(N2835), .B(N2905));
INVXL inst_cellmath__43_0_I390 (.Y(N2989), .A(N2835));
INVXL inst_cellmath__43_0_I391 (.Y(N3263), .A(a_man[4]));
NOR2XL inst_cellmath__43_0_I392 (.Y(N2666), .A(N3263), .B(N3303));
NOR2XL inst_cellmath__43_0_I393 (.Y(N1558), .A(N3263), .B(N1765));
NOR2XL inst_cellmath__43_0_I394 (.Y(N2417), .A(N3263), .B(N2196));
NOR2XL inst_cellmath__43_0_I395 (.Y(N3272), .A(N3263), .B(N2623));
NOR2XL inst_cellmath__43_0_I396 (.Y(N2165), .A(N3263), .B(N3050));
NOR2XL inst_cellmath__43_0_I397 (.Y(N3019), .A(N3263), .B(N3477));
NOR2XL inst_cellmath__43_0_I398 (.Y(N1913), .A(N3263), .B(N1948));
NOR2XL inst_cellmath__43_0_I399 (.Y(N2771), .A(N3263), .B(N2375));
NOR2XL inst_cellmath__43_0_I400 (.Y(N1666), .A(N3263), .B(N2806));
NOR2XL inst_cellmath__43_0_I401 (.Y(N2523), .A(N3263), .B(N3228));
NOR2XL inst_cellmath__43_0_I402 (.Y(N3376), .A(N3263), .B(N1702));
NOR2XL inst_cellmath__43_0_I403 (.Y(N2269), .A(N3263), .B(N2122));
NOR2XL inst_cellmath__43_0_I404 (.Y(N3124), .A(N3263), .B(N2556));
NOR2XL inst_cellmath__43_0_I405 (.Y(N2015), .A(N3263), .B(N2978));
NOR2XL inst_cellmath__43_0_I406 (.Y(N2875), .A(N3263), .B(N3412));
NOR2XL inst_cellmath__43_0_I407 (.Y(N1767), .A(N3263), .B(N1871));
NOR2XL inst_cellmath__43_0_I408 (.Y(N2625), .A(N3263), .B(N2301));
NOR2XL inst_cellmath__43_0_I409 (.Y(N3478), .A(N3263), .B(N2729));
NOR2XL inst_cellmath__43_0_I410 (.Y(N2378), .A(N3263), .B(N3157));
NOR2XL inst_cellmath__43_0_I411 (.Y(N3231), .A(N3263), .B(N1623));
NOR2XL inst_cellmath__43_0_I412 (.Y(N2123), .A(N3263), .B(N2049));
NOR2XL inst_cellmath__43_0_I413 (.Y(N2981), .A(N3263), .B(N2480));
NOR2XL inst_cellmath__43_0_I414 (.Y(N1874), .A(N3263), .B(N2905));
INVXL inst_cellmath__43_0_I415 (.Y(N2730), .A(N3263));
INVXL inst_cellmath__43_0_I416 (.Y(N1732), .A(a_man[5]));
NOR2XL inst_cellmath__43_0_I417 (.Y(N2409), .A(N1732), .B(N3303));
NOR2XL inst_cellmath__43_0_I418 (.Y(N3266), .A(N1732), .B(N1765));
NOR2XL inst_cellmath__43_0_I419 (.Y(N2158), .A(N1732), .B(N2196));
NOR2XL inst_cellmath__43_0_I420 (.Y(N3012), .A(N1732), .B(N2623));
NOR2XL inst_cellmath__43_0_I421 (.Y(N1907), .A(N1732), .B(N3050));
NOR2XL inst_cellmath__43_0_I422 (.Y(N2764), .A(N1732), .B(N3477));
NOR2XL inst_cellmath__43_0_I423 (.Y(N1659), .A(N1732), .B(N1948));
NOR2XL inst_cellmath__43_0_I424 (.Y(N2516), .A(N1732), .B(N2375));
NOR2XL inst_cellmath__43_0_I425 (.Y(N3369), .A(N1732), .B(N2806));
NOR2XL inst_cellmath__43_0_I426 (.Y(N2262), .A(N1732), .B(N3228));
NOR2XL inst_cellmath__43_0_I427 (.Y(N3116), .A(N1732), .B(N1702));
NOR2XL inst_cellmath__43_0_I428 (.Y(N2009), .A(N1732), .B(N2122));
NOR2XL inst_cellmath__43_0_I429 (.Y(N2867), .A(N1732), .B(N2556));
NOR2XL inst_cellmath__43_0_I430 (.Y(N1759), .A(N1732), .B(N2978));
NOR2XL inst_cellmath__43_0_I431 (.Y(N2617), .A(N1732), .B(N3412));
NOR2XL inst_cellmath__43_0_I432 (.Y(N3471), .A(N1732), .B(N1871));
NOR2XL inst_cellmath__43_0_I433 (.Y(N2369), .A(N1732), .B(N2301));
NOR2XL inst_cellmath__43_0_I434 (.Y(N3222), .A(N1732), .B(N2729));
NOR2XL inst_cellmath__43_0_I435 (.Y(N2114), .A(N1732), .B(N3157));
NOR2XL inst_cellmath__43_0_I436 (.Y(N2971), .A(N1732), .B(N1623));
NOR2XL inst_cellmath__43_0_I437 (.Y(N1865), .A(N1732), .B(N2049));
NOR2XL inst_cellmath__43_0_I438 (.Y(N2721), .A(N1732), .B(N2480));
NOR2XL inst_cellmath__43_0_I439 (.Y(N1618), .A(N1732), .B(N2905));
INVXL inst_cellmath__43_0_I440 (.Y(N2474), .A(N1732));
INVXL inst_cellmath__43_0_I441 (.Y(N2155), .A(a_man[6]));
NOR2XL inst_cellmath__43_0_I442 (.Y(N2148), .A(N2155), .B(N3303));
NOR2XL inst_cellmath__43_0_I443 (.Y(N3001), .A(N2155), .B(N1765));
NOR2XL inst_cellmath__43_0_I444 (.Y(N1894), .A(N2155), .B(N2196));
NOR2XL inst_cellmath__43_0_I445 (.Y(N2755), .A(N2155), .B(N2623));
NOR2XL inst_cellmath__43_0_I446 (.Y(N1648), .A(N2155), .B(N3050));
NOR2XL inst_cellmath__43_0_I447 (.Y(N2503), .A(N2155), .B(N3477));
NOR2XL inst_cellmath__43_0_I448 (.Y(N3361), .A(N2155), .B(N1948));
NOR2XL inst_cellmath__43_0_I449 (.Y(N2251), .A(N2155), .B(N2375));
NOR2XL inst_cellmath__43_0_I450 (.Y(N3105), .A(N2155), .B(N2806));
NOR2XL inst_cellmath__43_0_I451 (.Y(N2001), .A(N2155), .B(N3228));
NOR2XL inst_cellmath__43_0_I452 (.Y(N2857), .A(N2155), .B(N1702));
NOR2XL inst_cellmath__43_0_I453 (.Y(N1752), .A(N2155), .B(N2122));
NOR2XL inst_cellmath__43_0_I454 (.Y(N2608), .A(N2155), .B(N2556));
NOR2XL inst_cellmath__43_0_I455 (.Y(N3462), .A(N2155), .B(N2978));
NOR2XL inst_cellmath__43_0_I456 (.Y(N2361), .A(N2155), .B(N3412));
NOR2XL inst_cellmath__43_0_I457 (.Y(N3213), .A(N2155), .B(N1871));
NOR2XL inst_cellmath__43_0_I458 (.Y(N2106), .A(N2155), .B(N2301));
NOR2XL inst_cellmath__43_0_I459 (.Y(N2963), .A(N2155), .B(N2729));
NOR2XL inst_cellmath__43_0_I460 (.Y(N1856), .A(N2155), .B(N3157));
NOR2XL inst_cellmath__43_0_I461 (.Y(N2711), .A(N2155), .B(N1623));
NOR2XL inst_cellmath__43_0_I462 (.Y(N1609), .A(N2155), .B(N2049));
NOR2XL inst_cellmath__43_0_I463 (.Y(N2465), .A(N2155), .B(N2480));
NOR2XL inst_cellmath__43_0_I464 (.Y(N3318), .A(N2155), .B(N2905));
INVXL inst_cellmath__43_0_I465 (.Y(N2211), .A(N2155));
INVXL inst_cellmath__43_0_I466 (.Y(N2587), .A(a_man[7]));
NOR2XL inst_cellmath__43_0_I467 (.Y(N1886), .A(N2587), .B(N3303));
NOR2XL inst_cellmath__43_0_I468 (.Y(N2745), .A(N2587), .B(N1765));
NOR2XL inst_cellmath__43_0_I469 (.Y(N1640), .A(N2587), .B(N2196));
NOR2XL inst_cellmath__43_0_I470 (.Y(N2495), .A(N2587), .B(N2623));
NOR2XL inst_cellmath__43_0_I471 (.Y(N3351), .A(N2587), .B(N3050));
NOR2XL inst_cellmath__43_0_I472 (.Y(N2243), .A(N2587), .B(N3477));
NOR2XL inst_cellmath__43_0_I473 (.Y(N3096), .A(N2587), .B(N1948));
NOR2XL inst_cellmath__43_0_I474 (.Y(N1994), .A(N2587), .B(N2375));
NOR2XL inst_cellmath__43_0_I475 (.Y(N2850), .A(N2587), .B(N2806));
NOR2XL inst_cellmath__43_0_I476 (.Y(N1743), .A(N2587), .B(N3228));
NOR2XL inst_cellmath__43_0_I477 (.Y(N2601), .A(N2587), .B(N1702));
NOR2XL inst_cellmath__43_0_I478 (.Y(N3454), .A(N2587), .B(N2122));
NOR2XL inst_cellmath__43_0_I479 (.Y(N2350), .A(N2587), .B(N2556));
NOR2XL inst_cellmath__43_0_I480 (.Y(N3206), .A(N2587), .B(N2978));
NOR2XL inst_cellmath__43_0_I481 (.Y(N2098), .A(N2587), .B(N3412));
NOR2XL inst_cellmath__43_0_I482 (.Y(N2953), .A(N2587), .B(N1871));
NOR2XL inst_cellmath__43_0_I483 (.Y(N1849), .A(N2587), .B(N2301));
NOR2XL inst_cellmath__43_0_I484 (.Y(N2704), .A(N2587), .B(N2729));
NOR2XL inst_cellmath__43_0_I485 (.Y(N1602), .A(N2587), .B(N3157));
NOR2XL inst_cellmath__43_0_I486 (.Y(N2457), .A(N2587), .B(N1623));
NOR2XL inst_cellmath__43_0_I487 (.Y(N3310), .A(N2587), .B(N2049));
NOR2XL inst_cellmath__43_0_I488 (.Y(N2205), .A(N2587), .B(N2480));
NOR2XL inst_cellmath__43_0_I489 (.Y(N3059), .A(N2587), .B(N2905));
INVXL inst_cellmath__43_0_I490 (.Y(N1954), .A(N2587));
INVXL inst_cellmath__43_0_I491 (.Y(N3011), .A(a_man[8]));
NOR2XL inst_cellmath__43_0_I492 (.Y(N1631), .A(N3011), .B(N3303));
NOR2XL inst_cellmath__43_0_I493 (.Y(N2487), .A(N3011), .B(N1765));
NOR2XL inst_cellmath__43_0_I494 (.Y(N3343), .A(N3011), .B(N2196));
NOR2XL inst_cellmath__43_0_I495 (.Y(N2234), .A(N3011), .B(N2623));
NOR2XL inst_cellmath__43_0_I496 (.Y(N3088), .A(N3011), .B(N3050));
NOR2XL inst_cellmath__43_0_I497 (.Y(N1985), .A(N3011), .B(N3477));
NOR2XL inst_cellmath__43_0_I498 (.Y(N2841), .A(N3011), .B(N1948));
NOR2XL inst_cellmath__43_0_I499 (.Y(N1737), .A(N3011), .B(N2375));
NOR2XL inst_cellmath__43_0_I500 (.Y(N2593), .A(N3011), .B(N2806));
NOR2XL inst_cellmath__43_0_I501 (.Y(N3447), .A(N3011), .B(N3228));
NOR2XL inst_cellmath__43_0_I502 (.Y(N2341), .A(N3011), .B(N1702));
NOR2XL inst_cellmath__43_0_I503 (.Y(N3197), .A(N3011), .B(N2122));
NOR2XL inst_cellmath__43_0_I504 (.Y(N2089), .A(N3011), .B(N2556));
NOR2XL inst_cellmath__43_0_I505 (.Y(N2945), .A(N3011), .B(N2978));
NOR2XL inst_cellmath__43_0_I506 (.Y(N1841), .A(N3011), .B(N3412));
NOR2XL inst_cellmath__43_0_I507 (.Y(N2696), .A(N3011), .B(N1871));
NOR2XL inst_cellmath__43_0_I508 (.Y(N1591), .A(N3011), .B(N2301));
NOR2XL inst_cellmath__43_0_I509 (.Y(N2449), .A(N3011), .B(N2729));
NOR2XL inst_cellmath__43_0_I510 (.Y(N3302), .A(N3011), .B(N3157));
NOR2XL inst_cellmath__43_0_I511 (.Y(N2193), .A(N3011), .B(N1623));
NOR2XL inst_cellmath__43_0_I512 (.Y(N3049), .A(N3011), .B(N2049));
NOR2XL inst_cellmath__43_0_I513 (.Y(N1947), .A(N3011), .B(N2480));
NOR2XL inst_cellmath__43_0_I514 (.Y(N2803), .A(N3011), .B(N2905));
INVXL inst_cellmath__43_0_I515 (.Y(N1701), .A(N3011));
INVXL inst_cellmath__43_0_I516 (.Y(N3440), .A(a_man[9]));
NOR2XL inst_cellmath__43_0_I517 (.Y(N3334), .A(N3440), .B(N3303));
NOR2XL inst_cellmath__43_0_I518 (.Y(N2225), .A(N3440), .B(N1765));
NOR2XL inst_cellmath__43_0_I519 (.Y(N3080), .A(N3440), .B(N2196));
NOR2XL inst_cellmath__43_0_I520 (.Y(N1978), .A(N3440), .B(N2623));
NOR2XL inst_cellmath__43_0_I521 (.Y(N2834), .A(N3440), .B(N3050));
NOR2XL inst_cellmath__43_0_I522 (.Y(N1730), .A(N3440), .B(N3477));
NOR2XL inst_cellmath__43_0_I523 (.Y(N2586), .A(N3440), .B(N1948));
NOR2XL inst_cellmath__43_0_I524 (.Y(N3439), .A(N3440), .B(N2375));
NOR2XL inst_cellmath__43_0_I525 (.Y(N2333), .A(N3440), .B(N2806));
NOR2XL inst_cellmath__43_0_I526 (.Y(N3189), .A(N3440), .B(N3228));
NOR2XL inst_cellmath__43_0_I527 (.Y(N2080), .A(N3440), .B(N1702));
NOR2XL inst_cellmath__43_0_I528 (.Y(N2936), .A(N3440), .B(N2122));
NOR2XL inst_cellmath__43_0_I529 (.Y(N1832), .A(N3440), .B(N2556));
NOR2XL inst_cellmath__43_0_I530 (.Y(N2687), .A(N3440), .B(N2978));
NOR2XL inst_cellmath__43_0_I531 (.Y(N1582), .A(N3440), .B(N3412));
NOR2XL inst_cellmath__43_0_I532 (.Y(N2442), .A(N3440), .B(N1871));
NOR2XL inst_cellmath__43_0_I533 (.Y(N3293), .A(N3440), .B(N2301));
NOR2XL inst_cellmath__43_0_I534 (.Y(N2185), .A(N3440), .B(N2729));
NOR2XL inst_cellmath__43_0_I535 (.Y(N3041), .A(N3440), .B(N3157));
NOR2XL inst_cellmath__43_0_I536 (.Y(N1936), .A(N3440), .B(N1623));
NOR2XL inst_cellmath__43_0_I537 (.Y(N2794), .A(N3440), .B(N2049));
NOR2XL inst_cellmath__43_0_I538 (.Y(N1692), .A(N3440), .B(N2480));
NOR2XL inst_cellmath__43_0_I539 (.Y(N2547), .A(N3440), .B(N2905));
INVXL inst_cellmath__43_0_I540 (.Y(N3401), .A(N3440));
INVXL inst_cellmath__43_0_I541 (.Y(N1904), .A(a_man[10]));
NOR2XL inst_cellmath__43_0_I542 (.Y(N3071), .A(N1904), .B(N3303));
NOR2XL inst_cellmath__43_0_I543 (.Y(N1968), .A(N1904), .B(N1765));
NOR2XL inst_cellmath__43_0_I544 (.Y(N2825), .A(N1904), .B(N2196));
NOR2XL inst_cellmath__43_0_I545 (.Y(N1721), .A(N1904), .B(N2623));
NOR2XL inst_cellmath__43_0_I546 (.Y(N2577), .A(N1904), .B(N3050));
NOR2XL inst_cellmath__43_0_I547 (.Y(N3431), .A(N1904), .B(N3477));
NOR2XL inst_cellmath__43_0_I548 (.Y(N2324), .A(N1904), .B(N1948));
NOR2XL inst_cellmath__43_0_I549 (.Y(N3179), .A(N1904), .B(N2375));
NOR2XL inst_cellmath__43_0_I550 (.Y(N2070), .A(N1904), .B(N2806));
NOR2XL inst_cellmath__43_0_I551 (.Y(N2926), .A(N1904), .B(N3228));
NOR2XL inst_cellmath__43_0_I552 (.Y(N1822), .A(N1904), .B(N1702));
NOR2XL inst_cellmath__43_0_I553 (.Y(N2678), .A(N1904), .B(N2122));
NOR2XL inst_cellmath__43_0_I554 (.Y(N1571), .A(N1904), .B(N2556));
NOR2XL inst_cellmath__43_0_I555 (.Y(N2431), .A(N1904), .B(N2978));
NOR2XL inst_cellmath__43_0_I556 (.Y(N3283), .A(N1904), .B(N3412));
NOR2XL inst_cellmath__43_0_I557 (.Y(N2176), .A(N1904), .B(N1871));
NOR2XL inst_cellmath__43_0_I558 (.Y(N3031), .A(N1904), .B(N2301));
NOR2XL inst_cellmath__43_0_I559 (.Y(N1926), .A(N1904), .B(N2729));
NOR2XL inst_cellmath__43_0_I560 (.Y(N2784), .A(N1904), .B(N3157));
NOR2XL inst_cellmath__43_0_I561 (.Y(N1681), .A(N1904), .B(N1623));
NOR2XL inst_cellmath__43_0_I562 (.Y(N2537), .A(N1904), .B(N2049));
NOR2XL inst_cellmath__43_0_I563 (.Y(N3391), .A(N1904), .B(N2480));
NOR2XL inst_cellmath__43_0_I564 (.Y(N2283), .A(N1904), .B(N2905));
INVXL inst_cellmath__43_0_I565 (.Y(N3139), .A(N1904));
INVXL inst_cellmath__43_0_I566 (.Y(N2335), .A(a_man[11]));
NOR2XL inst_cellmath__43_0_I567 (.Y(N2817), .A(N2335), .B(N3303));
NOR2XL inst_cellmath__43_0_I568 (.Y(N1713), .A(N2335), .B(N1765));
NOR2XL inst_cellmath__43_0_I569 (.Y(N2568), .A(N2335), .B(N2196));
NOR2XL inst_cellmath__43_0_I570 (.Y(N3423), .A(N2335), .B(N2623));
NOR2XL inst_cellmath__43_0_I571 (.Y(N2315), .A(N2335), .B(N3050));
NOR2XL inst_cellmath__43_0_I572 (.Y(N3170), .A(N2335), .B(N3477));
NOR2XL inst_cellmath__43_0_I573 (.Y(N2062), .A(N2335), .B(N1948));
NOR2XL inst_cellmath__43_0_I574 (.Y(N2918), .A(N2335), .B(N2375));
NOR2XL inst_cellmath__43_0_I575 (.Y(N1812), .A(N2335), .B(N2806));
NOR2XL inst_cellmath__43_0_I576 (.Y(N2669), .A(N2335), .B(N3228));
NOR2XL inst_cellmath__43_0_I577 (.Y(N1561), .A(N2335), .B(N1702));
NOR2XL inst_cellmath__43_0_I578 (.Y(N2421), .A(N2335), .B(N2122));
NOR2XL inst_cellmath__43_0_I579 (.Y(N3275), .A(N2335), .B(N2556));
NOR2XL inst_cellmath__43_0_I580 (.Y(N2168), .A(N2335), .B(N2978));
NOR2XL inst_cellmath__43_0_I581 (.Y(N3023), .A(N2335), .B(N3412));
NOR2XL inst_cellmath__43_0_I582 (.Y(N1916), .A(N2335), .B(N1871));
NOR2XL inst_cellmath__43_0_I583 (.Y(N2774), .A(N2335), .B(N2301));
NOR2XL inst_cellmath__43_0_I584 (.Y(N1671), .A(N2335), .B(N2729));
NOR2XL inst_cellmath__43_0_I585 (.Y(N2527), .A(N2335), .B(N3157));
NOR2XL inst_cellmath__43_0_I586 (.Y(N3379), .A(N2335), .B(N1623));
NOR2XL inst_cellmath__43_0_I587 (.Y(N2274), .A(N2335), .B(N2049));
NOR2XL inst_cellmath__43_0_I588 (.Y(N3128), .A(N2335), .B(N2480));
NOR2XL inst_cellmath__43_0_I589 (.Y(N2018), .A(N2335), .B(N2905));
INVXL inst_cellmath__43_0_I590 (.Y(N2880), .A(N2335));
INVXL inst_cellmath__43_0_I591 (.Y(N2762), .A(a_man[12]));
NOR2XL inst_cellmath__43_0_I592 (.Y(N2561), .A(N2762), .B(N3303));
NOR2XL inst_cellmath__43_0_I593 (.Y(N3417), .A(N2762), .B(N1765));
NOR2XL inst_cellmath__43_0_I594 (.Y(N2305), .A(N2762), .B(N2196));
NOR2XL inst_cellmath__43_0_I595 (.Y(N3163), .A(N2762), .B(N2623));
NOR2XL inst_cellmath__43_0_I596 (.Y(N2055), .A(N2762), .B(N3050));
NOR2XL inst_cellmath__43_0_I597 (.Y(N2910), .A(N2762), .B(N3477));
NOR2XL inst_cellmath__43_0_I598 (.Y(N1805), .A(N2762), .B(N1948));
NOR2XL inst_cellmath__43_0_I599 (.Y(N2662), .A(N2762), .B(N2375));
NOR2XL inst_cellmath__43_0_I600 (.Y(N1554), .A(N2762), .B(N2806));
NOR2XL inst_cellmath__43_0_I601 (.Y(N2413), .A(N2762), .B(N3228));
NOR2XL inst_cellmath__43_0_I602 (.Y(N3268), .A(N2762), .B(N1702));
NOR2XL inst_cellmath__43_0_I603 (.Y(N2161), .A(N2762), .B(N2122));
NOR2XL inst_cellmath__43_0_I604 (.Y(N3015), .A(N2762), .B(N2556));
NOR2XL inst_cellmath__43_0_I605 (.Y(N1909), .A(N2762), .B(N2978));
NOR2XL inst_cellmath__43_0_I606 (.Y(N2767), .A(N2762), .B(N3412));
NOR2XL inst_cellmath__43_0_I607 (.Y(N1662), .A(N2762), .B(N1871));
NOR2XL inst_cellmath__43_0_I608 (.Y(N2519), .A(N2762), .B(N2301));
NOR2XL inst_cellmath__43_0_I609 (.Y(N3372), .A(N2762), .B(N2729));
NOR2XL inst_cellmath__43_0_I610 (.Y(N2265), .A(N2762), .B(N3157));
NOR2XL inst_cellmath__43_0_I611 (.Y(N3119), .A(N2762), .B(N1623));
NOR2XL inst_cellmath__43_0_I612 (.Y(N2012), .A(N2762), .B(N2049));
NOR2XL inst_cellmath__43_0_I613 (.Y(N2873), .A(N2762), .B(N2480));
NOR2XL inst_cellmath__43_0_I614 (.Y(N1762), .A(N2762), .B(N2905));
INVXL inst_cellmath__43_0_I615 (.Y(N2620), .A(N2762));
INVXL inst_cellmath__43_0_I616 (.Y(N3190), .A(a_man[13]));
NOR2XL inst_cellmath__43_0_I617 (.Y(N2295), .A(N3190), .B(N3303));
NOR2XL inst_cellmath__43_0_I618 (.Y(N3152), .A(N3190), .B(N1765));
NOR2XL inst_cellmath__43_0_I619 (.Y(N2044), .A(N3190), .B(N2196));
NOR2XL inst_cellmath__43_0_I620 (.Y(N2900), .A(N3190), .B(N2623));
NOR2XL inst_cellmath__43_0_I621 (.Y(N1793), .A(N3190), .B(N3050));
NOR2XL inst_cellmath__43_0_I622 (.Y(N2655), .A(N3190), .B(N3477));
NOR2XL inst_cellmath__43_0_I623 (.Y(N3507), .A(N3190), .B(N1948));
NOR2XL inst_cellmath__43_0_I624 (.Y(N2402), .A(N3190), .B(N2375));
NOR2XL inst_cellmath__43_0_I625 (.Y(N3259), .A(N3190), .B(N2806));
NOR2XL inst_cellmath__43_0_I626 (.Y(N2151), .A(N3190), .B(N3228));
NOR2XL inst_cellmath__43_0_I627 (.Y(N3005), .A(N3190), .B(N1702));
NOR2XL inst_cellmath__43_0_I628 (.Y(N1900), .A(N3190), .B(N2122));
NOR2XL inst_cellmath__43_0_I629 (.Y(N2758), .A(N3190), .B(N2556));
NOR2XL inst_cellmath__43_0_I630 (.Y(N1652), .A(N3190), .B(N2978));
NOR2XL inst_cellmath__43_0_I631 (.Y(N2509), .A(N3190), .B(N3412));
NOR2XL inst_cellmath__43_0_I632 (.Y(N3364), .A(N3190), .B(N1871));
NOR2XL inst_cellmath__43_0_I633 (.Y(N2255), .A(N3190), .B(N2301));
NOR2XL inst_cellmath__43_0_I634 (.Y(N3111), .A(N3190), .B(N2729));
NOR2XL inst_cellmath__43_0_I635 (.Y(N2005), .A(N3190), .B(N3157));
NOR2XL inst_cellmath__43_0_I636 (.Y(N2861), .A(N3190), .B(N1623));
NOR2XL inst_cellmath__43_0_I637 (.Y(N1755), .A(N3190), .B(N2049));
NOR2XL inst_cellmath__43_0_I638 (.Y(N2613), .A(N3190), .B(N2480));
NOR2XL inst_cellmath__43_0_I639 (.Y(N3466), .A(N3190), .B(N2905));
INVXL inst_cellmath__43_0_I640 (.Y(N2365), .A(N3190));
INVXL inst_cellmath__43_0_I641 (.Y(N1658), .A(a_man[14]));
NOR2XL inst_cellmath__43_0_I642 (.Y(N2036), .A(N1658), .B(N3303));
NOR2XL inst_cellmath__43_0_I643 (.Y(N2892), .A(N1658), .B(N1765));
NOR2XL inst_cellmath__43_0_I644 (.Y(N1783), .A(N1658), .B(N2196));
NOR2XL inst_cellmath__43_0_I645 (.Y(N2644), .A(N1658), .B(N2623));
NOR2XL inst_cellmath__43_0_I646 (.Y(N3497), .A(N1658), .B(N3050));
NOR2XL inst_cellmath__43_0_I647 (.Y(N2392), .A(N1658), .B(N3477));
NOR2XL inst_cellmath__43_0_I648 (.Y(N3250), .A(N1658), .B(N1948));
NOR2XL inst_cellmath__43_0_I649 (.Y(N2141), .A(N1658), .B(N2375));
NOR2XL inst_cellmath__43_0_I650 (.Y(N2996), .A(N1658), .B(N2806));
NOR2XL inst_cellmath__43_0_I651 (.Y(N1891), .A(N1658), .B(N3228));
NOR2XL inst_cellmath__43_0_I652 (.Y(N2748), .A(N1658), .B(N1702));
NOR2XL inst_cellmath__43_0_I653 (.Y(N1643), .A(N1658), .B(N2122));
NOR2XL inst_cellmath__43_0_I654 (.Y(N2500), .A(N1658), .B(N2556));
NOR2XL inst_cellmath__43_0_I655 (.Y(N3354), .A(N1658), .B(N2978));
NOR2XL inst_cellmath__43_0_I656 (.Y(N2246), .A(N1658), .B(N3412));
NOR2XL inst_cellmath__43_0_I657 (.Y(N3101), .A(N1658), .B(N1871));
NOR2XL inst_cellmath__43_0_I658 (.Y(N1997), .A(N1658), .B(N2301));
NOR2XL inst_cellmath__43_0_I659 (.Y(N2853), .A(N1658), .B(N2729));
NOR2XL inst_cellmath__43_0_I660 (.Y(N1747), .A(N1658), .B(N3157));
NOR2XL inst_cellmath__43_0_I661 (.Y(N2604), .A(N1658), .B(N1623));
NOR2XL inst_cellmath__43_0_I662 (.Y(N3457), .A(N1658), .B(N2049));
NOR2XL inst_cellmath__43_0_I663 (.Y(N2357), .A(N1658), .B(N2480));
NOR2XL inst_cellmath__43_0_I664 (.Y(N3209), .A(N1658), .B(N2905));
INVXL inst_cellmath__43_0_I665 (.Y(N2102), .A(N1658));
INVXL inst_cellmath__43_0_I666 (.Y(N2081), .A(a_man[15]));
NOR2XL inst_cellmath__43_0_I667 (.Y(N1775), .A(N2081), .B(N3303));
NOR2XL inst_cellmath__43_0_I668 (.Y(N2633), .A(N2081), .B(N1765));
NOR2XL inst_cellmath__43_0_I669 (.Y(N3489), .A(N2081), .B(N2196));
NOR2XL inst_cellmath__43_0_I670 (.Y(N2385), .A(N2081), .B(N2623));
NOR2XL inst_cellmath__43_0_I671 (.Y(N3238), .A(N2081), .B(N3050));
NOR2XL inst_cellmath__43_0_I672 (.Y(N2133), .A(N2081), .B(N3477));
NOR2XL inst_cellmath__43_0_I673 (.Y(N2988), .A(N2081), .B(N1948));
NOR2XL inst_cellmath__43_0_I674 (.Y(N1882), .A(N2081), .B(N2375));
NOR2XL inst_cellmath__43_0_I675 (.Y(N2740), .A(N2081), .B(N2806));
NOR2XL inst_cellmath__43_0_I676 (.Y(N1634), .A(N2081), .B(N3228));
NOR2XL inst_cellmath__43_0_I677 (.Y(N2492), .A(N2081), .B(N1702));
NOR2XL inst_cellmath__43_0_I678 (.Y(N3345), .A(N2081), .B(N2122));
NOR2XL inst_cellmath__43_0_I679 (.Y(N2236), .A(N2081), .B(N2556));
NOR2XL inst_cellmath__43_0_I680 (.Y(N3092), .A(N2081), .B(N2978));
NOR2XL inst_cellmath__43_0_I681 (.Y(N1987), .A(N2081), .B(N3412));
NOR2XL inst_cellmath__43_0_I682 (.Y(N2844), .A(N2081), .B(N1871));
NOR2XL inst_cellmath__43_0_I683 (.Y(N1741), .A(N2081), .B(N2301));
NOR2XL inst_cellmath__43_0_I684 (.Y(N2595), .A(N2081), .B(N2729));
NOR2XL inst_cellmath__43_0_I685 (.Y(N3449), .A(N2081), .B(N3157));
NOR2XL inst_cellmath__43_0_I686 (.Y(N2345), .A(N2081), .B(N1623));
NOR2XL inst_cellmath__43_0_I687 (.Y(N3199), .A(N2081), .B(N2049));
NOR2XL inst_cellmath__43_0_I688 (.Y(N2092), .A(N2081), .B(N2480));
NOR2XL inst_cellmath__43_0_I689 (.Y(N2949), .A(N2081), .B(N2905));
INVXL inst_cellmath__43_0_I690 (.Y(N1843), .A(N2081));
INVXL inst_cellmath__43_0_I691 (.Y(N2513), .A(a_man[16]));
NOR2XL inst_cellmath__43_0_I692 (.Y(N3481), .A(N2513), .B(N3303));
NOR2XL inst_cellmath__43_0_I693 (.Y(N2377), .A(N2513), .B(N1765));
NOR2XL inst_cellmath__43_0_I694 (.Y(N3230), .A(N2513), .B(N2196));
NOR2XL inst_cellmath__43_0_I695 (.Y(N2126), .A(N2513), .B(N2623));
NOR2XL inst_cellmath__43_0_I696 (.Y(N2980), .A(N2513), .B(N3050));
NOR2XL inst_cellmath__43_0_I697 (.Y(N1873), .A(N2513), .B(N3477));
NOR2XL inst_cellmath__43_0_I698 (.Y(N2733), .A(N2513), .B(N1948));
NOR2XL inst_cellmath__43_0_I699 (.Y(N1626), .A(N2513), .B(N2375));
NOR2XL inst_cellmath__43_0_I700 (.Y(N2482), .A(N2513), .B(N2806));
NOR2XL inst_cellmath__43_0_I701 (.Y(N3338), .A(N2513), .B(N3228));
NOR2XL inst_cellmath__43_0_I702 (.Y(N2229), .A(N2513), .B(N1702));
NOR2XL inst_cellmath__43_0_I703 (.Y(N3082), .A(N2513), .B(N2122));
NOR2XL inst_cellmath__43_0_I704 (.Y(N1981), .A(N2513), .B(N2556));
NOR2XL inst_cellmath__43_0_I705 (.Y(N2838), .A(N2513), .B(N2978));
NOR2XL inst_cellmath__43_0_I706 (.Y(N1733), .A(N2513), .B(N3412));
NOR2XL inst_cellmath__43_0_I707 (.Y(N2590), .A(N2513), .B(N1871));
NOR2XL inst_cellmath__43_0_I708 (.Y(N3442), .A(N2513), .B(N2301));
NOR2XL inst_cellmath__43_0_I709 (.Y(N2338), .A(N2513), .B(N2729));
NOR2XL inst_cellmath__43_0_I710 (.Y(N3192), .A(N2513), .B(N3157));
NOR2XL inst_cellmath__43_0_I711 (.Y(N2083), .A(N2513), .B(N1623));
NOR2XL inst_cellmath__43_0_I712 (.Y(N2941), .A(N2513), .B(N2049));
NOR2XL inst_cellmath__43_0_I713 (.Y(N1835), .A(N2513), .B(N2480));
NOR2XL inst_cellmath__43_0_I714 (.Y(N2690), .A(N2513), .B(N2905));
INVXL inst_cellmath__43_0_I715 (.Y(N1587), .A(N2513));
INVXL inst_cellmath__43_0_I716 (.Y(N2938), .A(a_man[17]));
NOR2XL inst_cellmath__43_0_I717 (.Y(N3221), .A(N2938), .B(N3303));
NOR2XL inst_cellmath__43_0_I718 (.Y(N2117), .A(N2938), .B(N1765));
NOR2XL inst_cellmath__43_0_I719 (.Y(N2970), .A(N2938), .B(N2196));
NOR2XL inst_cellmath__43_0_I720 (.Y(N1864), .A(N2938), .B(N2623));
NOR2XL inst_cellmath__43_0_I721 (.Y(N2724), .A(N2938), .B(N3050));
NOR2XL inst_cellmath__43_0_I722 (.Y(N1617), .A(N2938), .B(N3477));
NOR2XL inst_cellmath__43_0_I723 (.Y(N2473), .A(N2938), .B(N1948));
NOR2XL inst_cellmath__43_0_I724 (.Y(N3329), .A(N2938), .B(N2375));
NOR2XL inst_cellmath__43_0_I725 (.Y(N2220), .A(N2938), .B(N2806));
NOR2XL inst_cellmath__43_0_I726 (.Y(N3073), .A(N2938), .B(N3228));
NOR2XL inst_cellmath__43_0_I727 (.Y(N1973), .A(N2938), .B(N1702));
NOR2XL inst_cellmath__43_0_I728 (.Y(N2828), .A(N2938), .B(N2122));
NOR2XL inst_cellmath__43_0_I729 (.Y(N1723), .A(N2938), .B(N2556));
NOR2XL inst_cellmath__43_0_I730 (.Y(N2581), .A(N2938), .B(N2978));
NOR2XL inst_cellmath__43_0_I731 (.Y(N3434), .A(N2938), .B(N3412));
NOR2XL inst_cellmath__43_0_I732 (.Y(N2326), .A(N2938), .B(N1871));
NOR2XL inst_cellmath__43_0_I733 (.Y(N3183), .A(N2938), .B(N2301));
NOR2XL inst_cellmath__43_0_I734 (.Y(N2074), .A(N2938), .B(N2729));
NOR2XL inst_cellmath__43_0_I735 (.Y(N2928), .A(N2938), .B(N3157));
NOR2XL inst_cellmath__43_0_I736 (.Y(N1826), .A(N2938), .B(N1623));
NOR2XL inst_cellmath__43_0_I737 (.Y(N2681), .A(N2938), .B(N2049));
NOR2XL inst_cellmath__43_0_I738 (.Y(N1574), .A(N2938), .B(N2480));
NOR2XL inst_cellmath__43_0_I739 (.Y(N2436), .A(N2938), .B(N2905));
INVXL inst_cellmath__43_0_I740 (.Y(N3286), .A(N2938));
INVXL inst_cellmath__43_0_I741 (.Y(N3367), .A(a_man[18]));
NOR2XL inst_cellmath__43_0_I742 (.Y(N2962), .A(N3367), .B(N3303));
NOR2XL inst_cellmath__43_0_I743 (.Y(N1855), .A(N3367), .B(N1765));
NOR2XL inst_cellmath__43_0_I744 (.Y(N2714), .A(N3367), .B(N2196));
NOR2XL inst_cellmath__43_0_I745 (.Y(N1608), .A(N3367), .B(N2623));
NOR2XL inst_cellmath__43_0_I746 (.Y(N2464), .A(N3367), .B(N3050));
NOR2XL inst_cellmath__43_0_I747 (.Y(N3321), .A(N3367), .B(N3477));
NOR2XL inst_cellmath__43_0_I748 (.Y(N2210), .A(N3367), .B(N1948));
NOR2XL inst_cellmath__43_0_I749 (.Y(N3065), .A(N3367), .B(N2375));
NOR2XL inst_cellmath__43_0_I750 (.Y(N1964), .A(N3367), .B(N2806));
NOR2XL inst_cellmath__43_0_I751 (.Y(N2819), .A(N3367), .B(N3228));
NOR2XL inst_cellmath__43_0_I752 (.Y(N1715), .A(N3367), .B(N1702));
NOR2XL inst_cellmath__43_0_I753 (.Y(N2572), .A(N3367), .B(N2122));
NOR2XL inst_cellmath__43_0_I754 (.Y(N3425), .A(N3367), .B(N2556));
NOR2XL inst_cellmath__43_0_I755 (.Y(N2318), .A(N3367), .B(N2978));
NOR2XL inst_cellmath__43_0_I756 (.Y(N3174), .A(N3367), .B(N3412));
NOR2XL inst_cellmath__43_0_I757 (.Y(N2065), .A(N3367), .B(N1871));
NOR2XL inst_cellmath__43_0_I758 (.Y(N2920), .A(N3367), .B(N2301));
NOR2XL inst_cellmath__43_0_I759 (.Y(N1816), .A(N3367), .B(N2729));
NOR2XL inst_cellmath__43_0_I760 (.Y(N2672), .A(N3367), .B(N3157));
NOR2XL inst_cellmath__43_0_I761 (.Y(N1564), .A(N3367), .B(N1623));
NOR2XL inst_cellmath__43_0_I762 (.Y(N2426), .A(N3367), .B(N2049));
NOR2XL inst_cellmath__43_0_I763 (.Y(N3277), .A(N3367), .B(N2480));
NOR2XL inst_cellmath__43_0_I764 (.Y(N2170), .A(N3367), .B(N2905));
INVXL inst_cellmath__43_0_I765 (.Y(N3026), .A(N3367));
INVXL inst_cellmath__43_0_I766 (.Y(N1833), .A(a_man[19]));
NOR2XL inst_cellmath__43_0_I767 (.Y(N2703), .A(N1833), .B(N3303));
NOR2XL inst_cellmath__43_0_I768 (.Y(N1601), .A(N1833), .B(N1765));
NOR2XL inst_cellmath__43_0_I769 (.Y(N2456), .A(N1833), .B(N2196));
NOR2XL inst_cellmath__43_0_I770 (.Y(N3314), .A(N1833), .B(N2623));
NOR2XL inst_cellmath__43_0_I771 (.Y(N2204), .A(N1833), .B(N3050));
NOR2XL inst_cellmath__43_0_I772 (.Y(N3058), .A(N1833), .B(N3477));
NOR2XL inst_cellmath__43_0_I773 (.Y(N1957), .A(N1833), .B(N1948));
NOR2XL inst_cellmath__43_0_I774 (.Y(N2813), .A(N1833), .B(N2375));
NOR2XL inst_cellmath__43_0_I775 (.Y(N1708), .A(N1833), .B(N2806));
NOR2XL inst_cellmath__43_0_I776 (.Y(N2565), .A(N1833), .B(N3228));
NOR2XL inst_cellmath__43_0_I777 (.Y(N3419), .A(N1833), .B(N1702));
NOR2XL inst_cellmath__43_0_I778 (.Y(N2309), .A(N1833), .B(N2122));
NOR2XL inst_cellmath__43_0_I779 (.Y(N3167), .A(N1833), .B(N2556));
NOR2XL inst_cellmath__43_0_I780 (.Y(N2057), .A(N1833), .B(N2978));
NOR2XL inst_cellmath__43_0_I781 (.Y(N2914), .A(N1833), .B(N3412));
NOR2XL inst_cellmath__43_0_I782 (.Y(N1809), .A(N1833), .B(N1871));
NOR2XL inst_cellmath__43_0_I783 (.Y(N2664), .A(N1833), .B(N2301));
NOR2XL inst_cellmath__43_0_I784 (.Y(N1556), .A(N1833), .B(N2729));
NOR2XL inst_cellmath__43_0_I785 (.Y(N2416), .A(N1833), .B(N3157));
NOR2XL inst_cellmath__43_0_I786 (.Y(N3270), .A(N1833), .B(N1623));
NOR2XL inst_cellmath__43_0_I787 (.Y(N2163), .A(N1833), .B(N2049));
NOR2XL inst_cellmath__43_0_I788 (.Y(N3018), .A(N1833), .B(N2480));
NOR2XL inst_cellmath__43_0_I789 (.Y(N1911), .A(N1833), .B(N2905));
INVXL inst_cellmath__43_0_I790 (.Y(N2769), .A(N1833));
INVXL inst_cellmath__43_0_I791 (.Y(N2261), .A(a_man[20]));
NOR2XL inst_cellmath__43_0_I792 (.Y(N2448), .A(N2261), .B(N3303));
NOR2XL inst_cellmath__43_0_I793 (.Y(N3301), .A(N2261), .B(N1765));
NOR2XL inst_cellmath__43_0_I794 (.Y(N2195), .A(N2261), .B(N2196));
NOR2XL inst_cellmath__43_0_I795 (.Y(N3048), .A(N2261), .B(N2623));
NOR2XL inst_cellmath__43_0_I796 (.Y(N1946), .A(N2261), .B(N3050));
NOR2XL inst_cellmath__43_0_I797 (.Y(N2805), .A(N2261), .B(N3477));
NOR2XL inst_cellmath__43_0_I798 (.Y(N1700), .A(N2261), .B(N1948));
NOR2XL inst_cellmath__43_0_I799 (.Y(N2555), .A(N2261), .B(N2375));
NOR2XL inst_cellmath__43_0_I800 (.Y(N3411), .A(N2261), .B(N2806));
NOR2XL inst_cellmath__43_0_I801 (.Y(N2300), .A(N2261), .B(N3228));
NOR2XL inst_cellmath__43_0_I802 (.Y(N3159), .A(N2261), .B(N1702));
NOR2XL inst_cellmath__43_0_I803 (.Y(N2048), .A(N2261), .B(N2122));
NOR2XL inst_cellmath__43_0_I804 (.Y(N2904), .A(N2261), .B(N2556));
NOR2XL inst_cellmath__43_0_I805 (.Y(N1801), .A(N2261), .B(N2978));
NOR2XL inst_cellmath__43_0_I806 (.Y(N2658), .A(N2261), .B(N3412));
NOR2XL inst_cellmath__43_0_I807 (.Y(N3511), .A(N2261), .B(N1871));
NOR2XL inst_cellmath__43_0_I808 (.Y(N2407), .A(N2261), .B(N2301));
NOR2XL inst_cellmath__43_0_I809 (.Y(N3262), .A(N2261), .B(N2729));
NOR2XL inst_cellmath__43_0_I810 (.Y(N2154), .A(N2261), .B(N3157));
NOR2XL inst_cellmath__43_0_I811 (.Y(N3010), .A(N2261), .B(N1623));
NOR2XL inst_cellmath__43_0_I812 (.Y(N1903), .A(N2261), .B(N2049));
NOR2XL inst_cellmath__43_0_I813 (.Y(N2761), .A(N2261), .B(N2480));
NOR2XL inst_cellmath__43_0_I814 (.Y(N1657), .A(N2261), .B(N2905));
INVXL inst_cellmath__43_0_I815 (.Y(N2512), .A(N2261));
INVXL inst_cellmath__43_0_I816 (.Y(N2688), .A(a_man[21]));
NOR2XL inst_cellmath__43_0_I817 (.Y(N2187), .A(N2688), .B(N3303));
NOR2XL inst_cellmath__43_0_I818 (.Y(N3040), .A(N2688), .B(N1765));
NOR2XL inst_cellmath__43_0_I819 (.Y(N1935), .A(N2688), .B(N2196));
NOR2XL inst_cellmath__43_0_I820 (.Y(N2796), .A(N2688), .B(N2623));
NOR2XL inst_cellmath__43_0_I821 (.Y(N1691), .A(N2688), .B(N3050));
NOR2XL inst_cellmath__43_0_I822 (.Y(N2546), .A(N2688), .B(N3477));
NOR2XL inst_cellmath__43_0_I823 (.Y(N3403), .A(N2688), .B(N1948));
NOR2XL inst_cellmath__43_0_I824 (.Y(N2291), .A(N2688), .B(N2375));
NOR2XL inst_cellmath__43_0_I825 (.Y(N3147), .A(N2688), .B(N2806));
NOR2XL inst_cellmath__43_0_I826 (.Y(N2038), .A(N2688), .B(N3228));
NOR2XL inst_cellmath__43_0_I827 (.Y(N2896), .A(N2688), .B(N1702));
NOR2XL inst_cellmath__43_0_I828 (.Y(N1787), .A(N2688), .B(N2122));
NOR2XL inst_cellmath__43_0_I829 (.Y(N2648), .A(N2688), .B(N2556));
NOR2XL inst_cellmath__43_0_I830 (.Y(N3502), .A(N2688), .B(N2978));
NOR2XL inst_cellmath__43_0_I831 (.Y(N2397), .A(N2688), .B(N3412));
NOR2XL inst_cellmath__43_0_I832 (.Y(N3253), .A(N2688), .B(N1871));
NOR2XL inst_cellmath__43_0_I833 (.Y(N2145), .A(N2688), .B(N2301));
NOR2XL inst_cellmath__43_0_I834 (.Y(N2999), .A(N2688), .B(N2729));
NOR2XL inst_cellmath__43_0_I835 (.Y(N1893), .A(N2688), .B(N3157));
NOR2XL inst_cellmath__43_0_I836 (.Y(N2751), .A(N2688), .B(N1623));
NOR2XL inst_cellmath__43_0_I837 (.Y(N1647), .A(N2688), .B(N2049));
NOR2XL inst_cellmath__43_0_I838 (.Y(N2502), .A(N2688), .B(N2480));
NOR2XL inst_cellmath__43_0_I839 (.Y(N3357), .A(N2688), .B(N2905));
INVXL inst_cellmath__43_0_I840 (.Y(N2250), .A(N2688));
INVXL inst_cellmath__43_0_I841 (.Y(N3114), .A(a_man[22]));
NOR2XL inst_cellmath__43_0_I842 (.Y(N1925), .A(N3114), .B(N3303));
NOR2XL inst_cellmath__43_0_I843 (.Y(N2786), .A(N3114), .B(N1765));
NOR2XL inst_cellmath__43_0_I844 (.Y(N1680), .A(N3114), .B(N2196));
NOR2XL inst_cellmath__43_0_I845 (.Y(N2536), .A(N3114), .B(N2623));
NOR2XL inst_cellmath__43_0_I846 (.Y(N3393), .A(N3114), .B(N3050));
NOR2XL inst_cellmath__43_0_I847 (.Y(N2282), .A(N3114), .B(N3477));
NOR2XL inst_cellmath__43_0_I848 (.Y(N3138), .A(N3114), .B(N1948));
NOR2XL inst_cellmath__43_0_I849 (.Y(N2029), .A(N3114), .B(N2375));
NOR2XL inst_cellmath__43_0_I850 (.Y(N2888), .A(N3114), .B(N2806));
NOR2XL inst_cellmath__43_0_I851 (.Y(N1779), .A(N3114), .B(N3228));
NOR2XL inst_cellmath__43_0_I852 (.Y(N2638), .A(N3114), .B(N1702));
NOR2XL inst_cellmath__43_0_I853 (.Y(N3492), .A(N3114), .B(N2122));
NOR2XL inst_cellmath__43_0_I854 (.Y(N2388), .A(N3114), .B(N2556));
NOR2XL inst_cellmath__43_0_I855 (.Y(N3244), .A(N3114), .B(N2978));
NOR2XL inst_cellmath__43_0_I856 (.Y(N2137), .A(N3114), .B(N3412));
NOR2XL inst_cellmath__43_0_I857 (.Y(N2991), .A(N3114), .B(N1871));
NOR2XL inst_cellmath__43_0_I858 (.Y(N1885), .A(N3114), .B(N2301));
NOR2XL inst_cellmath__43_0_I859 (.Y(N2743), .A(N3114), .B(N2729));
NOR2XL inst_cellmath__43_0_I860 (.Y(N1638), .A(N3114), .B(N3157));
NOR2XL inst_cellmath__43_0_I861 (.Y(N2494), .A(N3114), .B(N1623));
NOR2XL inst_cellmath__43_0_I862 (.Y(N3349), .A(N3114), .B(N2049));
NOR2XL inst_cellmath__43_0_I863 (.Y(N2240), .A(N3114), .B(N2480));
NOR2XL inst_cellmath__43_0_I864 (.Y(N3094), .A(N3114), .B(N2905));
INVXL inst_cellmath__43_0_I865 (.Y(N1991), .A(N3114));
INVXL inst_cellmath__43_0_I866 (.Y(N1915), .A(N3303));
INVXL inst_cellmath__43_0_I867 (.Y(N2776), .A(N1765));
INVXL inst_cellmath__43_0_I868 (.Y(N1670), .A(N2196));
INVXL inst_cellmath__43_0_I869 (.Y(N2526), .A(N2623));
INVXL inst_cellmath__43_0_I870 (.Y(N3381), .A(N3050));
INVXL inst_cellmath__43_0_I871 (.Y(N2273), .A(N3477));
INVXL inst_cellmath__43_0_I872 (.Y(N3127), .A(N1948));
INVXL inst_cellmath__43_0_I873 (.Y(N2020), .A(N2375));
INVXL inst_cellmath__43_0_I874 (.Y(N2879), .A(N2806));
INVXL inst_cellmath__43_0_I875 (.Y(N1769), .A(N3228));
INVXL inst_cellmath__43_0_I876 (.Y(N2629), .A(N1702));
INVXL inst_cellmath__43_0_I877 (.Y(N3483), .A(N2122));
INVXL inst_cellmath__43_0_I878 (.Y(N2380), .A(N2556));
INVXL inst_cellmath__43_0_I879 (.Y(N3235), .A(N2978));
INVXL inst_cellmath__43_0_I880 (.Y(N2128), .A(N3412));
INVXL inst_cellmath__43_0_I881 (.Y(N2983), .A(N1871));
INVXL inst_cellmath__43_0_I882 (.Y(N1878), .A(N2301));
INVXL inst_cellmath__43_0_I883 (.Y(N2736), .A(N2729));
INVXL inst_cellmath__43_0_I884 (.Y(N1628), .A(N3157));
INVXL inst_cellmath__43_0_I885 (.Y(N2486), .A(N1623));
INVXL inst_cellmath__43_0_I886 (.Y(N3341), .A(N2049));
INVXL inst_cellmath__43_0_I887 (.Y(N2231), .A(N2480));
INVXL inst_cellmath__43_0_I888 (.Y(N3087), .A(N2905));
ADDHX1 inst_cellmath__43_0_I889 (.CO(N2371), .S(N1945), .A(N3452), .B(N2339));
ADDHX1 inst_cellmath__43_0_I890 (.CO(N3227), .S(N2801), .A(N2347), .B(N3194));
ADDFX1 inst_cellmath__43_0_I891 (.CO(N2119), .S(N1695), .A(N2077), .B(N2923), .CI(N2371));
ADDHX1 inst_cellmath__43_0_I892 (.CO(N2973), .S(N2554), .A(N3201), .B(N2086));
ADDFX1 inst_cellmath__43_0_I893 (.CO(N1870), .S(N3408), .A(N1817), .B(N2932), .CI(N2666));
ADDFX1 inst_cellmath__43_0_I894 (.CO(N2726), .S(N2294), .A(N2554), .B(N3227), .CI(N2119));
ADDHX1 inst_cellmath__43_0_I895 (.CO(N1620), .S(N3156), .A(N2096), .B(N2942));
ADDFX1 inst_cellmath__43_0_I896 (.CO(N2479), .S(N2043), .A(N2675), .B(N1827), .CI(N1558));
ADDFX1 inst_cellmath__43_0_I897 (.CO(N3331), .S(N2899), .A(N2973), .B(N2409), .CI(N3156));
ADDFX1 inst_cellmath__43_0_I898 (.CO(N2222), .S(N1797), .A(N2043), .B(N1870), .CI(N2899));
ADDHX1 inst_cellmath__43_0_I899 (.CO(N3079), .S(N2654), .A(N2951), .B(N1837));
ADDFX1 inst_cellmath__43_0_I900 (.CO(N1975), .S(N3506), .A(N1567), .B(N2685), .CI(N2417));
ADDFX1 inst_cellmath__43_0_I901 (.CO(N2830), .S(N2405), .A(N2148), .B(N3266), .CI(N1620));
ADDFX1 inst_cellmath__43_0_I902 (.CO(N1729), .S(N3258), .A(N2479), .B(N2654), .CI(N3506));
ADDFX1 inst_cellmath__43_0_I903 (.CO(N2583), .S(N2150), .A(N2405), .B(N3331), .CI(N3258));
ADDHX1 inst_cellmath__43_0_I904 (.CO(N3436), .S(N3008), .A(N1845), .B(N2693));
ADDFX1 inst_cellmath__43_0_I905 (.CO(N2332), .S(N1899), .A(N2427), .B(N1578), .CI(N3272));
ADDFX1 inst_cellmath__43_0_I906 (.CO(N3186), .S(N2757), .A(N3001), .B(N2158), .CI(N1886));
ADDFX1 inst_cellmath__43_0_I907 (.CO(N2076), .S(N1655), .A(N3008), .B(N3079), .CI(N1975));
ADDFX1 inst_cellmath__43_0_I908 (.CO(N2935), .S(N2508), .A(N1899), .B(N2830), .CI(N2757));
ADDFX1 inst_cellmath__43_0_I909 (.CO(N1829), .S(N3363), .A(N1655), .B(N1729), .CI(N2508));
ADDHX1 inst_cellmath__43_0_I910 (.CO(N2684), .S(N2258), .A(N2701), .B(N1588));
ADDFX1 inst_cellmath__43_0_I911 (.CO(N1581), .S(N3110), .A(N3280), .B(N2437), .CI(N2165));
ADDFX1 inst_cellmath__43_0_I912 (.CO(N2439), .S(N2004), .A(N1894), .B(N3012), .CI(N2745));
ADDFX1 inst_cellmath__43_0_I913 (.CO(N3289), .S(N2864), .A(N3436), .B(N1631), .CI(N2258));
ADDFX1 inst_cellmath__43_0_I914 (.CO(N2184), .S(N1754), .A(N3186), .B(N2332), .CI(N3110));
ADDFX1 inst_cellmath__43_0_I915 (.CO(N3037), .S(N2612), .A(N2076), .B(N2004), .CI(N2864));
ADDFX1 inst_cellmath__43_0_I916 (.CO(N1931), .S(N3469), .A(N1754), .B(N2935), .CI(N2612));
ADDHX1 inst_cellmath__43_0_I917 (.CO(N2793), .S(N2364), .A(N1596), .B(N2446));
ADDFX1 inst_cellmath__43_0_I918 (.CO(N1687), .S(N3217), .A(N2173), .B(N3290), .CI(N3019));
ADDFX1 inst_cellmath__43_0_I919 (.CO(N2542), .S(N2112), .A(N2755), .B(N1907), .CI(N1640));
ADDFX1 inst_cellmath__43_0_I920 (.CO(N3400), .S(N2966), .A(N3334), .B(N2487), .CI(N2684));
ADDFX1 inst_cellmath__43_0_I921 (.CO(N2287), .S(N1860), .A(N1581), .B(N2364), .CI(N2439));
ADDFX1 inst_cellmath__43_0_I922 (.CO(N3143), .S(N2717), .A(N2112), .B(N3217), .CI(N3289));
ADDFX1 inst_cellmath__43_0_I923 (.CO(N2035), .S(N1612), .A(N2184), .B(N2966), .CI(N1860));
ADDFX1 inst_cellmath__43_0_I924 (.CO(N2891), .S(N2470), .A(N3037), .B(N2717), .CI(N1612));
ADDHX1 inst_cellmath__43_0_I925 (.CO(N1786), .S(N3324), .A(N2452), .B(N3298));
ADDFX1 inst_cellmath__43_0_I926 (.CO(N2643), .S(N2213), .A(N3027), .B(N2181), .CI(N1913));
ADDFX1 inst_cellmath__43_0_I927 (.CO(N3496), .S(N3070), .A(N1648), .B(N2764), .CI(N2495));
ADDFX1 inst_cellmath__43_0_I928 (.CO(N2396), .S(N1966), .A(N2225), .B(N3343), .CI(N3071));
ADDFX1 inst_cellmath__43_0_I929 (.CO(N3249), .S(N2821), .A(N3324), .B(N2793), .CI(N1687));
ADDFX1 inst_cellmath__43_0_I930 (.CO(N2140), .S(N1720), .A(N3400), .B(N2542), .CI(N2213));
ADDFX1 inst_cellmath__43_0_I931 (.CO(N2998), .S(N2575), .A(N1966), .B(N3070), .CI(N2287));
ADDFX1 inst_cellmath__43_0_I932 (.CO(N1890), .S(N3427), .A(N3143), .B(N2821), .CI(N1720));
ADDFX1 inst_cellmath__43_0_I933 (.CO(N2747), .S(N2323), .A(N2035), .B(N2575), .CI(N3427));
ADDHX1 inst_cellmath__43_0_I934 (.CO(N1645), .S(N3176), .A(N3308), .B(N2190));
ADDFX1 inst_cellmath__43_0_I935 (.CO(N2499), .S(N2067), .A(N1922), .B(N3035), .CI(N2771));
ADDFX1 inst_cellmath__43_0_I936 (.CO(N3353), .S(N2925), .A(N2503), .B(N1659), .CI(N3351));
ADDFX1 inst_cellmath__43_0_I937 (.CO(N2248), .S(N1819), .A(N3080), .B(N2234), .CI(N1968));
ADDFX1 inst_cellmath__43_0_I938 (.CO(N3100), .S(N2674), .A(N1786), .B(N2817), .CI(N3176));
ADDFX1 inst_cellmath__43_0_I939 (.CO(N1996), .S(N1570), .A(N3496), .B(N2643), .CI(N2396));
ADDFX1 inst_cellmath__43_0_I940 (.CO(N2855), .S(N2429), .A(N2925), .B(N2067), .CI(N1819));
ADDFX1 inst_cellmath__43_0_I941 (.CO(N1746), .S(N3279), .A(N2674), .B(N3249), .CI(N2140));
ADDFX1 inst_cellmath__43_0_I942 (.CO(N2603), .S(N2175), .A(N2998), .B(N1570), .CI(N2429));
ADDFX1 inst_cellmath__43_0_I943 (.CO(N3460), .S(N3029), .A(N1890), .B(N3279), .CI(N2175));
ADDHX1 inst_cellmath__43_0_I944 (.CO(N2356), .S(N1921), .A(N2199), .B(N3044));
ADDFX1 inst_cellmath__43_0_I945 (.CO(N3208), .S(N2783), .A(N2780), .B(N1932), .CI(N1666));
ADDFX1 inst_cellmath__43_0_I946 (.CO(N2104), .S(N1677), .A(N3361), .B(N2516), .CI(N2243));
ADDFX1 inst_cellmath__43_0_I947 (.CO(N2958), .S(N2533), .A(N1978), .B(N3088), .CI(N2825));
ADDFX1 inst_cellmath__43_0_I948 (.CO(N1852), .S(N3390), .A(N2561), .B(N1713), .CI(N1645));
ADDFX1 inst_cellmath__43_0_I949 (.CO(N2709), .S(N2280), .A(N2499), .B(N1921), .CI(N3353));
ADDFX1 inst_cellmath__43_0_I950 (.CO(N1604), .S(N3134), .A(N2783), .B(N2248), .CI(N1677));
ADDFX1 inst_cellmath__43_0_I951 (.CO(N2460), .S(N2027), .A(N3100), .B(N2533), .CI(N3390));
ADDFX1 inst_cellmath__43_0_I952 (.CO(N3316), .S(N2886), .A(N2855), .B(N1996), .CI(N2280));
ADDFX1 inst_cellmath__43_0_I953 (.CO(N2207), .S(N1774), .A(N1746), .B(N3134), .CI(N2027));
ADDFX1 inst_cellmath__43_0_I954 (.CO(N3062), .S(N2636), .A(N2886), .B(N2603), .CI(N1774));
ADDHX1 inst_cellmath__43_0_I955 (.CO(N1959), .S(N3488), .A(N3055), .B(N1942));
ADDFX1 inst_cellmath__43_0_I956 (.CO(N2815), .S(N2384), .A(N1675), .B(N2790), .CI(N2523));
ADDFX1 inst_cellmath__43_0_I957 (.CO(N1710), .S(N3242), .A(N2251), .B(N3369), .CI(N3096));
ADDFX1 inst_cellmath__43_0_I958 (.CO(N2567), .S(N2132), .A(N2834), .B(N1985), .CI(N1721));
ADDFX1 inst_cellmath__43_0_I959 (.CO(N3421), .S(N2987), .A(N3417), .B(N2568), .CI(N2295));
ADDFX1 inst_cellmath__43_0_I960 (.CO(N2311), .S(N1881), .A(N3488), .B(N2356), .CI(N3208));
ADDFX1 inst_cellmath__43_0_I961 (.CO(N3169), .S(N2739), .A(N2958), .B(N2104), .CI(N1852));
ADDFX1 inst_cellmath__43_0_I962 (.CO(N2058), .S(N1637), .A(N3242), .B(N2384), .CI(N2132));
ADDFX1 inst_cellmath__43_0_I963 (.CO(N2917), .S(N2491), .A(N2709), .B(N2987), .CI(N1881));
ADDFX1 inst_cellmath__43_0_I964 (.CO(N1811), .S(N3344), .A(N2460), .B(N1604), .CI(N2739));
ADDFX1 inst_cellmath__43_0_I965 (.CO(N2665), .S(N2239), .A(N3316), .B(N1637), .CI(N2491));
ADDFX1 inst_cellmath__43_0_I966 (.CO(N1560), .S(N3091), .A(N2207), .B(N3344), .CI(N2239));
ADDHX1 inst_cellmath__43_0_I967 (.CO(N2419), .S(N1986), .A(N1952), .B(N2799));
ADDFX1 inst_cellmath__43_0_I968 (.CO(N3271), .S(N2847), .A(N2534), .B(N1685), .CI(N3376));
ADDFX1 inst_cellmath__43_0_I969 (.CO(N2167), .S(N1740), .A(N3105), .B(N2262), .CI(N1994));
ADDFX1 inst_cellmath__43_0_I970 (.CO(N3021), .S(N2594), .A(N1730), .B(N2841), .CI(N2577));
ADDFX1 inst_cellmath__43_0_I971 (.CO(N1912), .S(N3451), .A(N2305), .B(N3423), .CI(N3152));
ADDFX1 inst_cellmath__43_0_I972 (.CO(N2773), .S(N2344), .A(N1959), .B(N2036), .CI(N1986));
ADDFX1 inst_cellmath__43_0_I973 (.CO(N1668), .S(N3198), .A(N1710), .B(N2815), .CI(N2567));
ADDFX1 inst_cellmath__43_0_I974 (.CO(N2522), .S(N2095), .A(N2847), .B(N3421), .CI(N1740));
ADDFX1 inst_cellmath__43_0_I975 (.CO(N3378), .S(N2948), .A(N3451), .B(N2594), .CI(N2311));
ADDFX1 inst_cellmath__43_0_I976 (.CO(N2271), .S(N1842), .A(N3169), .B(N2344), .CI(N2058));
ADDFX1 inst_cellmath__43_0_I977 (.CO(N3122), .S(N2700), .A(N2095), .B(N3198), .CI(N2948));
ADDFX1 inst_cellmath__43_0_I978 (.CO(N2017), .S(N1594), .A(N1811), .B(N2917), .CI(N1842));
ADDFX1 inst_cellmath__43_0_I979 (.CO(N2877), .S(N2450), .A(N2665), .B(N2700), .CI(N1594));
ADDHX1 inst_cellmath__43_0_I980 (.CO(N1766), .S(N3307), .A(N2810), .B(N1696));
ADDFX1 inst_cellmath__43_0_I981 (.CO(N2627), .S(N2198), .A(N3387), .B(N2543), .CI(N2269));
ADDFX1 inst_cellmath__43_0_I982 (.CO(N3480), .S(N3052), .A(N2001), .B(N3116), .CI(N2850));
ADDFX1 inst_cellmath__43_0_I983 (.CO(N2376), .S(N1951), .A(N2586), .B(N1737), .CI(N3431));
ADDFX1 inst_cellmath__43_0_I984 (.CO(N3233), .S(N2808), .A(N3163), .B(N2315), .CI(N2044));
ADDFX1 inst_cellmath__43_0_I985 (.CO(N2125), .S(N1703), .A(N1775), .B(N2892), .CI(N2419));
ADDFX1 inst_cellmath__43_0_I986 (.CO(N2979), .S(N2560), .A(N3271), .B(N3307), .CI(N2167));
ADDFX1 inst_cellmath__43_0_I987 (.CO(N1876), .S(N3414), .A(N1912), .B(N3021), .CI(N2198));
ADDFX1 inst_cellmath__43_0_I988 (.CO(N2732), .S(N2302), .A(N1951), .B(N3052), .CI(N2808));
ADDFX1 inst_cellmath__43_0_I989 (.CO(N1625), .S(N3162), .A(N1703), .B(N2773), .CI(N1668));
ADDFX1 inst_cellmath__43_0_I990 (.CO(N2484), .S(N2052), .A(N2560), .B(N2522), .CI(N3378));
ADDFX1 inst_cellmath__43_0_I991 (.CO(N3337), .S(N2907), .A(N2302), .B(N3414), .CI(N2271));
ADDFX1 inst_cellmath__43_0_I992 (.CO(N2228), .S(N1804), .A(N2052), .B(N3162), .CI(N3122));
ADDFX1 inst_cellmath__43_0_I993 (.CO(N3084), .S(N2660), .A(N2017), .B(N2907), .CI(N1804));
ADDHX1 inst_cellmath__43_0_I994 (.CO(N1980), .S(N1551), .A(N1705), .B(N2551));
ADDFX1 inst_cellmath__43_0_I995 (.CO(N2837), .S(N2412), .A(N2278), .B(N3397), .CI(N3124));
ADDFX1 inst_cellmath__43_0_I996 (.CO(N1735), .S(N3265), .A(N2857), .B(N2009), .CI(N1743));
ADDFX1 inst_cellmath__43_0_I997 (.CO(N2589), .S(N2157), .A(N3439), .B(N2593), .CI(N2324));
ADDFX1 inst_cellmath__43_0_I998 (.CO(N3444), .S(N3014), .A(N2055), .B(N3170), .CI(N2900));
ADDFX1 inst_cellmath__43_0_I999 (.CO(N2337), .S(N1906), .A(N2633), .B(N1783), .CI(N3481));
ADDFX1 inst_cellmath__43_0_I1000 (.CO(N3191), .S(N2766), .A(N1551), .B(N1766), .CI(N2627));
ADDFX1 inst_cellmath__43_0_I1001 (.CO(N2085), .S(N1661), .A(N2376), .B(N3480), .CI(N3233));
ADDFX1 inst_cellmath__43_0_I1002 (.CO(N2940), .S(N2515), .A(N2412), .B(N2125), .CI(N3265));
ADDFX1 inst_cellmath__43_0_I1003 (.CO(N1834), .S(N3371), .A(N3014), .B(N2157), .CI(N1906));
ADDFX1 inst_cellmath__43_0_I1004 (.CO(N2692), .S(N2264), .A(N1876), .B(N2979), .CI(N2732));
ADDFX1 inst_cellmath__43_0_I1005 (.CO(N1586), .S(N3115), .A(N1661), .B(N2766), .CI(N1625));
ADDFX1 inst_cellmath__43_0_I1006 (.CO(N2443), .S(N2011), .A(N3371), .B(N2515), .CI(N2484));
ADDFX1 inst_cellmath__43_0_I1007 (.CO(N3297), .S(N2869), .A(N3337), .B(N2264), .CI(N3115));
ADDFX1 inst_cellmath__43_0_I1008 (.CO(N2189), .S(N1758), .A(N2228), .B(N2011), .CI(N2869));
ADDHX1 inst_cellmath__43_0_I1009 (.CO(N3042), .S(N2619), .A(N2562), .B(N3406));
ADDFX1 inst_cellmath__43_0_I1010 (.CO(N1940), .S(N3473), .A(N3135), .B(N2288), .CI(N2015));
ADDFX1 inst_cellmath__43_0_I1011 (.CO(N2798), .S(N2368), .A(N1752), .B(N2867), .CI(N2601));
ADDFX1 inst_cellmath__43_0_I1012 (.CO(N1693), .S(N3224), .A(N2333), .B(N3447), .CI(N3179));
ADDFX1 inst_cellmath__43_0_I1013 (.CO(N2550), .S(N2116), .A(N2910), .B(N2062), .CI(N1793));
ADDFX1 inst_cellmath__43_0_I1014 (.CO(N3405), .S(N2969), .A(N3489), .B(N2644), .CI(N2377));
ADDFX1 inst_cellmath__43_0_I1015 (.CO(N2292), .S(N1867), .A(N1980), .B(N3221), .CI(N2619));
ADDFX1 inst_cellmath__43_0_I1016 (.CO(N3151), .S(N2723), .A(N1735), .B(N2837), .CI(N2589));
ADDFX1 inst_cellmath__43_0_I1017 (.CO(N2040), .S(N1616), .A(N2337), .B(N3444), .CI(N3473));
ADDFX1 inst_cellmath__43_0_I1018 (.CO(N2897), .S(N2476), .A(N3224), .B(N2368), .CI(N2116));
ADDFX1 inst_cellmath__43_0_I1019 (.CO(N1792), .S(N3328), .A(N3191), .B(N2969), .CI(N2085));
ADDFX1 inst_cellmath__43_0_I1020 (.CO(N2651), .S(N2219), .A(N2940), .B(N1867), .CI(N2723));
ADDFX1 inst_cellmath__43_0_I1021 (.CO(N3504), .S(N3076), .A(N1616), .B(N1834), .CI(N2476));
ADDFX1 inst_cellmath__43_0_I1022 (.CO(N2401), .S(N1972), .A(N3328), .B(N2692), .CI(N1586));
ADDFX1 inst_cellmath__43_0_I1023 (.CO(N3256), .S(N2827), .A(N3076), .B(N2219), .CI(N2443));
ADDFX1 inst_cellmath__43_0_I1024 (.CO(N2147), .S(N1726), .A(N3297), .B(N1972), .CI(N2827));
ADDHX1 inst_cellmath__43_0_I1025 (.CO(N3004), .S(N2580), .A(N3415), .B(N2296));
ADDFX1 inst_cellmath__43_0_I1026 (.CO(N1897), .S(N3433), .A(N2024), .B(N3144), .CI(N2875));
ADDFX1 inst_cellmath__43_0_I1027 (.CO(N2754), .S(N2329), .A(N2608), .B(N1759), .CI(N3454));
ADDFX1 inst_cellmath__43_0_I1028 (.CO(N1651), .S(N3182), .A(N3189), .B(N2341), .CI(N2070));
ADDFX1 inst_cellmath__43_0_I1029 (.CO(N2506), .S(N2073), .A(N1805), .B(N2918), .CI(N2655));
ADDFX1 inst_cellmath__43_0_I1030 (.CO(N3360), .S(N2931), .A(N2385), .B(N3497), .CI(N3230));
ADDFX1 inst_cellmath__43_0_I1031 (.CO(N2254), .S(N1825), .A(N2962), .B(N2117), .CI(N3042));
ADDFX1 inst_cellmath__43_0_I1032 (.CO(N3108), .S(N2680), .A(N1940), .B(N2580), .CI(N2798));
ADDFX1 inst_cellmath__43_0_I1033 (.CO(N2000), .S(N1577), .A(N2550), .B(N1693), .CI(N3405));
ADDFX1 inst_cellmath__43_0_I1034 (.CO(N2860), .S(N2435), .A(N2329), .B(N3433), .CI(N3182));
ADDFX1 inst_cellmath__43_0_I1035 (.CO(N1751), .S(N3285), .A(N2931), .B(N2073), .CI(N2292));
ADDFX1 inst_cellmath__43_0_I1036 (.CO(N2611), .S(N2180), .A(N3151), .B(N1825), .CI(N2040));
ADDFX1 inst_cellmath__43_0_I1037 (.CO(N3465), .S(N3034), .A(N2680), .B(N2897), .CI(N1577));
ADDFX1 inst_cellmath__43_0_I1038 (.CO(N2360), .S(N1930), .A(N2435), .B(N1792), .CI(N3285));
ADDFX1 inst_cellmath__43_0_I1039 (.CO(N3216), .S(N2789), .A(N2180), .B(N2651), .CI(N3504));
ADDFX1 inst_cellmath__43_0_I1040 (.CO(N2109), .S(N1683), .A(N1930), .B(N3034), .CI(N2401));
ADDFX1 inst_cellmath__43_0_I1041 (.CO(N2961), .S(N2541), .A(N3256), .B(N2789), .CI(N1683));
ADDHX1 inst_cellmath__43_0_I1042 (.CO(N1859), .S(N3396), .A(N2306), .B(N3153));
ADDFX1 inst_cellmath__43_0_I1043 (.CO(N2713), .S(N2284), .A(N2884), .B(N2032), .CI(N1767));
ADDFX1 inst_cellmath__43_0_I1044 (.CO(N1607), .S(N3142), .A(N3462), .B(N2617), .CI(N2350));
ADDFX1 inst_cellmath__43_0_I1045 (.CO(N2467), .S(N2031), .A(N2080), .B(N3197), .CI(N2926));
ADDFX1 inst_cellmath__43_0_I1046 (.CO(N3320), .S(N2889), .A(N2662), .B(N1812), .CI(N3507));
ADDFX1 inst_cellmath__43_0_I1047 (.CO(N2209), .S(N1782), .A(N3238), .B(N2392), .CI(N2126));
ADDFX1 inst_cellmath__43_0_I1048 (.CO(N3067), .S(N2640), .A(N1855), .B(N2970), .CI(N2703));
ADDFX1 inst_cellmath__43_0_I1049 (.CO(N1963), .S(N3493), .A(N3396), .B(N3004), .CI(N1897));
ADDFX1 inst_cellmath__43_0_I1050 (.CO(N2818), .S(N2391), .A(N1651), .B(N2754), .CI(N2506));
ADDFX1 inst_cellmath__43_0_I1051 (.CO(N1717), .S(N3246), .A(N2254), .B(N3360), .CI(N2284));
ADDFX1 inst_cellmath__43_0_I1052 (.CO(N2571), .S(N2138), .A(N2031), .B(N3142), .CI(N2889));
ADDFX1 inst_cellmath__43_0_I1053 (.CO(N3424), .S(N2995), .A(N2640), .B(N1782), .CI(N3108));
ADDFX1 inst_cellmath__43_0_I1054 (.CO(N2320), .S(N1888), .A(N3493), .B(N2000), .CI(N2860));
ADDFX1 inst_cellmath__43_0_I1055 (.CO(N3173), .S(N2744), .A(N1751), .B(N2391), .CI(N3246));
ADDFX1 inst_cellmath__43_0_I1056 (.CO(N2064), .S(N1642), .A(N2611), .B(N2138), .CI(N2995));
ADDFX1 inst_cellmath__43_0_I1057 (.CO(N2922), .S(N2497), .A(N1888), .B(N3465), .CI(N2360));
ADDFX1 inst_cellmath__43_0_I1058 (.CO(N1815), .S(N3350), .A(N1642), .B(N2744), .CI(N3216));
ADDFX1 inst_cellmath__43_0_I1059 (.CO(N2671), .S(N2245), .A(N2109), .B(N2497), .CI(N3350));
ADDHX1 inst_cellmath__43_0_I1060 (.CO(N1566), .S(N3098), .A(N3164), .B(N2041));
ADDFX1 inst_cellmath__43_0_I1061 (.CO(N2425), .S(N1993), .A(N1776), .B(N2893), .CI(N2625));
ADDFX1 inst_cellmath__43_0_I1062 (.CO(N3276), .S(N2852), .A(N2361), .B(N3471), .CI(N3206));
ADDFX1 inst_cellmath__43_0_I1063 (.CO(N2172), .S(N1744), .A(N2936), .B(N2089), .CI(N1822));
ADDFX1 inst_cellmath__43_0_I1064 (.CO(N3025), .S(N2600), .A(N1554), .B(N2669), .CI(N2402));
ADDFX1 inst_cellmath__43_0_I1065 (.CO(N1919), .S(N3456), .A(N2133), .B(N3250), .CI(N2980));
ADDFX1 inst_cellmath__43_0_I1066 (.CO(N2779), .S(N2353), .A(N2714), .B(N1864), .CI(N1601));
ADDFX1 inst_cellmath__43_0_I1067 (.CO(N1674), .S(N3205), .A(N1859), .B(N2448), .CI(N3098));
ADDFX1 inst_cellmath__43_0_I1068 (.CO(N2531), .S(N2101), .A(N1607), .B(N2713), .CI(N2467));
ADDFX1 inst_cellmath__43_0_I1069 (.CO(N3385), .S(N2956), .A(N2209), .B(N3320), .CI(N3067));
ADDFX1 inst_cellmath__43_0_I1070 (.CO(N2277), .S(N1848), .A(N2852), .B(N1993), .CI(N1744));
ADDFX1 inst_cellmath__43_0_I1071 (.CO(N3131), .S(N2707), .A(N3456), .B(N2600), .CI(N2353));
ADDFX1 inst_cellmath__43_0_I1072 (.CO(N2023), .S(N1600), .A(N2818), .B(N1963), .CI(N3205));
ADDFX1 inst_cellmath__43_0_I1073 (.CO(N2883), .S(N2455), .A(N2101), .B(N1717), .CI(N2956));
ADDFX1 inst_cellmath__43_0_I1074 (.CO(N1773), .S(N3313), .A(N3424), .B(N2571), .CI(N1848));
ADDFX1 inst_cellmath__43_0_I1075 (.CO(N2632), .S(N2203), .A(N2320), .B(N2707), .CI(N1600));
ADDFX1 inst_cellmath__43_0_I1076 (.CO(N3485), .S(N3061), .A(N2455), .B(N3173), .CI(N2064));
ADDFX1 inst_cellmath__43_0_I1077 (.CO(N2383), .S(N1956), .A(N2922), .B(N3313), .CI(N2203));
ADDFX1 inst_cellmath__43_0_I1078 (.CO(N3237), .S(N2812), .A(N1815), .B(N3061), .CI(N1956));
ADDHX1 inst_cellmath__43_0_I1079 (.CO(N2129), .S(N1709), .A(N2053), .B(N2901));
ADDFX1 inst_cellmath__43_0_I1080 (.CO(N2986), .S(N2564), .A(N2634), .B(N1784), .CI(N3478));
ADDFX1 inst_cellmath__43_0_I1081 (.CO(N1879), .S(N3418), .A(N3213), .B(N2369), .CI(N2098));
ADDFX1 inst_cellmath__43_0_I1082 (.CO(N2737), .S(N2310), .A(N1832), .B(N2945), .CI(N2678));
ADDFX1 inst_cellmath__43_0_I1083 (.CO(N1633), .S(N3166), .A(N2413), .B(N1561), .CI(N3259));
ADDFX1 inst_cellmath__43_0_I1084 (.CO(N2488), .S(N2056), .A(N2988), .B(N2141), .CI(N1873));
ADDFX1 inst_cellmath__43_0_I1085 (.CO(N3342), .S(N2915), .A(N1608), .B(N2724), .CI(N2456));
ADDFX1 inst_cellmath__43_0_I1086 (.CO(N2235), .S(N1808), .A(N2187), .B(N3301), .CI(N1566));
ADDFX1 inst_cellmath__43_0_I1087 (.CO(N3089), .S(N2663), .A(N2425), .B(N1709), .CI(N3276));
ADDFX1 inst_cellmath__43_0_I1088 (.CO(N1984), .S(N1557), .A(N3025), .B(N2172), .CI(N1919));
ADDFX1 inst_cellmath__43_0_I1089 (.CO(N2843), .S(N2415), .A(N2564), .B(N2779), .CI(N3418));
ADDFX1 inst_cellmath__43_0_I1090 (.CO(N1738), .S(N3269), .A(N3166), .B(N2310), .CI(N2056));
ADDFX1 inst_cellmath__43_0_I1091 (.CO(N2592), .S(N2164), .A(N1674), .B(N2915), .CI(N1808));
ADDFX1 inst_cellmath__43_0_I1092 (.CO(N3448), .S(N3017), .A(N3385), .B(N2531), .CI(N2277));
ADDFX1 inst_cellmath__43_0_I1093 (.CO(N2342), .S(N1910), .A(N2663), .B(N3131), .CI(N1557));
ADDFX1 inst_cellmath__43_0_I1094 (.CO(N3196), .S(N2770), .A(N3269), .B(N2415), .CI(N2023));
ADDFX1 inst_cellmath__43_0_I1095 (.CO(N2091), .S(N1665), .A(N2883), .B(N2164), .CI(N3017));
ADDFX1 inst_cellmath__43_0_I1096 (.CO(N2946), .S(N2521), .A(N1910), .B(N1773), .CI(N2632));
ADDFX1 inst_cellmath__43_0_I1097 (.CO(N1840), .S(N3375), .A(N3485), .B(N2770), .CI(N1665));
ADDFX1 inst_cellmath__43_0_I1098 (.CO(N2697), .S(N2268), .A(N2383), .B(N2521), .CI(N3375));
XNOR2X1 inst_cellmath__43_0_I1099 (.Y(N3121), .A(N2911), .B(N1794));
OR2XL inst_cellmath__43_0_I1100 (.Y(N1592), .A(N2911), .B(N1794));
ADDFX1 inst_cellmath__43_0_I1101 (.CO(N3304), .S(N2874), .A(N3486), .B(N2641), .CI(N2378));
ADDFX1 inst_cellmath__43_0_I1102 (.CO(N2194), .S(N1764), .A(N2106), .B(N3222), .CI(N2953));
ADDFX1 inst_cellmath__43_0_I1103 (.CO(N3047), .S(N2624), .A(N2687), .B(N1841), .CI(N1571));
ADDFX1 inst_cellmath__43_0_I1104 (.CO(N1949), .S(N3476), .A(N3268), .B(N2421), .CI(N2151));
ADDFX1 inst_cellmath__43_0_I1105 (.CO(N2804), .S(N2374), .A(N1882), .B(N2996), .CI(N2733));
ADDFX1 inst_cellmath__43_0_I1106 (.CO(N1699), .S(N3229), .A(N2464), .B(N1617), .CI(N3314));
ADDFX1 inst_cellmath__43_0_I1107 (.CO(N2557), .S(N2121), .A(N3040), .B(N2195), .CI(N1925));
ADDFX1 inst_cellmath__43_0_I1108 (.CO(N3410), .S(N2976), .A(N3121), .B(N2129), .CI(N2986));
ADDFX1 inst_cellmath__43_0_I1109 (.CO(N2299), .S(N1872), .A(N2737), .B(N1879), .CI(N1633));
ADDFX1 inst_cellmath__43_0_I1110 (.CO(N3158), .S(N2728), .A(N3342), .B(N2488), .CI(N2235));
ADDFX1 inst_cellmath__43_0_I1111 (.CO(N2047), .S(N1624), .A(N1764), .B(N2874), .CI(N2624));
ADDFX1 inst_cellmath__43_0_I1112 (.CO(N2906), .S(N2481), .A(N2374), .B(N3476), .CI(N3229));
ADDFX1 inst_cellmath__43_0_I1113 (.CO(N1800), .S(N3333), .A(N3089), .B(N2121), .CI(N1984));
ADDFX1 inst_cellmath__43_0_I1114 (.CO(N2657), .S(N2227), .A(N2843), .B(N2976), .CI(N1872));
ADDFX1 inst_cellmath__43_0_I1115 (.CO(N3512), .S(N3081), .A(N2592), .B(N1738), .CI(N2728));
ADDFX1 inst_cellmath__43_0_I1116 (.CO(N2406), .S(N1977), .A(N2481), .B(N1624), .CI(N3448));
ADDFX1 inst_cellmath__43_0_I1117 (.CO(N3261), .S(N2836), .A(N3333), .B(N2342), .CI(N2227));
ADDFX1 inst_cellmath__43_0_I1118 (.CO(N2156), .S(N1731), .A(N3081), .B(N3196), .CI(N1977));
ADDFX1 inst_cellmath__43_0_I1119 (.CO(N3009), .S(N2585), .A(N2836), .B(N2091), .CI(N2946));
ADDFX1 inst_cellmath__43_0_I1120 (.CO(N1902), .S(N3441), .A(N1840), .B(N1731), .CI(N2585));
ADDHX1 inst_cellmath__43_0_I1121 (.CO(N2763), .S(N2334), .A(N1915), .B(N2652));
ADDFX1 inst_cellmath__43_0_I1122 (.CO(N1656), .S(N3188), .A(N3498), .B(N1806), .CI(N2386));
ADDFX1 inst_cellmath__43_0_I1123 (.CO(N2511), .S(N2082), .A(N2114), .B(N3231), .CI(N2963));
ADDFX1 inst_cellmath__43_0_I1124 (.CO(N3368), .S(N2937), .A(N2696), .B(N1849), .CI(N1582));
ADDFX1 inst_cellmath__43_0_I1125 (.CO(N2260), .S(N1830), .A(N3275), .B(N2431), .CI(N2161));
ADDFX1 inst_cellmath__43_0_I1126 (.CO(N3113), .S(N2689), .A(N1891), .B(N3005), .CI(N2740));
ADDFX1 inst_cellmath__43_0_I1127 (.CO(N2008), .S(N1583), .A(N2473), .B(N1626), .CI(N3321));
ADDFX1 inst_cellmath__43_0_I1128 (.CO(N2865), .S(N2441), .A(N3048), .B(N2204), .CI(N1935));
ADDFX1 inst_cellmath__43_0_I1129 (.CO(N1757), .S(N3295), .A(N1592), .B(N2786), .CI(N2334));
ADDFX1 inst_cellmath__43_0_I1130 (.CO(N2616), .S(N2186), .A(N2194), .B(N3304), .CI(N3047));
ADDFX1 inst_cellmath__43_0_I1131 (.CO(N3470), .S(N3039), .A(N2804), .B(N1949), .CI(N1699));
ADDFX1 inst_cellmath__43_0_I1132 (.CO(N2367), .S(N1938), .A(N3188), .B(N2557), .CI(N2082));
ADDFX1 inst_cellmath__43_0_I1133 (.CO(N3220), .S(N2795), .A(N1830), .B(N2937), .CI(N2689));
ADDFX1 inst_cellmath__43_0_I1134 (.CO(N2113), .S(N1690), .A(N2441), .B(N1583), .CI(N3410));
ADDFX1 inst_cellmath__43_0_I1135 (.CO(N2968), .S(N2548), .A(N3295), .B(N2299), .CI(N3158));
ADDFX1 inst_cellmath__43_0_I1136 (.CO(N1863), .S(N3402), .A(N2186), .B(N2047), .CI(N3039));
ADDFX1 inst_cellmath__43_0_I1137 (.CO(N2719), .S(N2290), .A(N1938), .B(N2906), .CI(N2795));
ADDFX1 inst_cellmath__43_0_I1138 (.CO(N1614), .S(N3149), .A(N1690), .B(N1800), .CI(N2657));
ADDFX1 inst_cellmath__43_0_I1139 (.CO(N2472), .S(N2037), .A(N3512), .B(N2548), .CI(N3402));
ADDFX1 inst_cellmath__43_0_I1140 (.CO(N3325), .S(N2895), .A(N2290), .B(N2406), .CI(N3149));
ADDFX1 inst_cellmath__43_0_I1141 (.CO(N2216), .S(N1788), .A(N2037), .B(N3261), .CI(N2156));
ADDFX1 inst_cellmath__43_0_I1142 (.CO(N3072), .S(N2647), .A(N3009), .B(N2895), .CI(N1788));
ADDHX1 inst_cellmath__43_0_I1143 (.CO(N1969), .S(N3501), .A(N2776), .B(N2393));
ADDFX1 inst_cellmath__43_0_I1144 (.CO(N2824), .S(N2398), .A(N3239), .B(N3508), .CI(N2123));
ADDFX1 inst_cellmath__43_0_I1145 (.CO(N1722), .S(N3252), .A(N1856), .B(N2971), .CI(N2704));
ADDFX1 inst_cellmath__43_0_I1146 (.CO(N2576), .S(N2144), .A(N2442), .B(N1591), .CI(N3283));
ADDFX1 inst_cellmath__43_0_I1147 (.CO(N3430), .S(N3000), .A(N3015), .B(N2168), .CI(N1900));
ADDFX1 inst_cellmath__43_0_I1148 (.CO(N2325), .S(N1892), .A(N1634), .B(N2748), .CI(N2482));
ADDFX1 inst_cellmath__43_0_I1149 (.CO(N3178), .S(N2752), .A(N2210), .B(N3329), .CI(N3058));
ADDFX1 inst_cellmath__43_0_I1150 (.CO(N2071), .S(N1646), .A(N2796), .B(N1946), .CI(N1680));
ADDFX1 inst_cellmath__43_0_I1151 (.CO(N2927), .S(N2501), .A(N3501), .B(N2763), .CI(N1656));
ADDFX1 inst_cellmath__43_0_I1152 (.CO(N1821), .S(N3358), .A(N3368), .B(N2511), .CI(N2260));
ADDFX1 inst_cellmath__43_0_I1153 (.CO(N2679), .S(N2249), .A(N2008), .B(N3113), .CI(N2865));
ADDFX1 inst_cellmath__43_0_I1154 (.CO(N1572), .S(N3103), .A(N3252), .B(N2398), .CI(N2144));
ADDFX1 inst_cellmath__43_0_I1155 (.CO(N2430), .S(N1999), .A(N1892), .B(N3000), .CI(N2752));
ADDFX1 inst_cellmath__43_0_I1156 (.CO(N3284), .S(N2856), .A(N1757), .B(N1646), .CI(N2616));
ADDFX1 inst_cellmath__43_0_I1157 (.CO(N2177), .S(N1748), .A(N2501), .B(N3470), .CI(N2367));
ADDFX1 inst_cellmath__43_0_I1158 (.CO(N3030), .S(N2606), .A(N3358), .B(N3220), .CI(N2249));
ADDFX1 inst_cellmath__43_0_I1159 (.CO(N1927), .S(N3461), .A(N3103), .B(N2113), .CI(N1999));
ADDFX1 inst_cellmath__43_0_I1160 (.CO(N2785), .S(N2358), .A(N2856), .B(N2968), .CI(N1863));
ADDFX1 inst_cellmath__43_0_I1161 (.CO(N1679), .S(N3212), .A(N2606), .B(N1748), .CI(N2719));
ADDFX1 inst_cellmath__43_0_I1162 (.CO(N2538), .S(N2105), .A(N3461), .B(N1614), .CI(N2472));
ADDFX1 inst_cellmath__43_0_I1163 (.CO(N3392), .S(N2959), .A(N3212), .B(N2358), .CI(N3325));
ADDFX1 inst_cellmath__43_0_I1164 (.CO(N2281), .S(N1854), .A(N2216), .B(N2105), .CI(N2959));
ADDFX1 inst_cellmath__43_0_I1165 (.CO(N3140), .S(N2710), .A(N2134), .B(N1670), .CI(N2981));
ADDFX1 inst_cellmath__43_0_I1166 (.CO(N2028), .S(N1606), .A(N1865), .B(N3247), .CI(N2711));
ADDFX1 inst_cellmath__43_0_I1167 (.CO(N2887), .S(N2463), .A(N2449), .B(N1602), .CI(N3293));
ADDFX1 inst_cellmath__43_0_I1168 (.CO(N1780), .S(N3317), .A(N3023), .B(N2176), .CI(N1909));
ADDFX1 inst_cellmath__43_0_I1169 (.CO(N2637), .S(N2208), .A(N1643), .B(N2758), .CI(N2492));
ADDFX1 inst_cellmath__43_0_I1170 (.CO(N3491), .S(N3064), .A(N2220), .B(N3338), .CI(N3065));
ADDFX1 inst_cellmath__43_0_I1171 (.CO(N2389), .S(N1960), .A(N2805), .B(N1957), .CI(N1691));
ADDFX1 inst_cellmath__43_0_I1172 (.CO(N3243), .S(N2816), .A(N1969), .B(N2536), .CI(N2824));
ADDFX1 inst_cellmath__43_0_I1173 (.CO(N2136), .S(N1714), .A(N2576), .B(N1722), .CI(N3430));
ADDFX1 inst_cellmath__43_0_I1174 (.CO(N2993), .S(N2569), .A(N3178), .B(N2325), .CI(N2071));
ADDFX1 inst_cellmath__43_0_I1175 (.CO(N1884), .S(N3422), .A(N1606), .B(N2710), .CI(N2463));
ADDFX1 inst_cellmath__43_0_I1176 (.CO(N2742), .S(N2317), .A(N2208), .B(N3317), .CI(N3064));
ADDFX1 inst_cellmath__43_0_I1177 (.CO(N1639), .S(N3171), .A(N2927), .B(N1960), .CI(N1821));
ADDFX1 inst_cellmath__43_0_I1178 (.CO(N2493), .S(N2061), .A(N2816), .B(N2679), .CI(N1572));
ADDFX1 inst_cellmath__43_0_I1179 (.CO(N3348), .S(N2919), .A(N1714), .B(N2430), .CI(N2569));
ADDFX1 inst_cellmath__43_0_I1180 (.CO(N2242), .S(N1813), .A(N3422), .B(N3284), .CI(N2317));
ADDFX1 inst_cellmath__43_0_I1181 (.CO(N3093), .S(N2668), .A(N3171), .B(N2177), .CI(N3030));
ADDFX1 inst_cellmath__43_0_I1182 (.CO(N1990), .S(N1563), .A(N2919), .B(N2061), .CI(N1927));
ADDFX1 inst_cellmath__43_0_I1183 (.CO(N2849), .S(N2422), .A(N1813), .B(N2785), .CI(N2668));
ADDFX1 inst_cellmath__43_0_I1184 (.CO(N1742), .S(N3274), .A(N1563), .B(N1679), .CI(N2538));
ADDFX1 inst_cellmath__43_0_I1185 (.CO(N2598), .S(N2169), .A(N3392), .B(N2422), .CI(N3274));
ADDFX1 inst_cellmath__43_0_I1186 (.CO(N3453), .S(N3022), .A(N1874), .B(N2526), .CI(N2721));
ADDFX1 inst_cellmath__43_0_I1187 (.CO(N2348), .S(N1918), .A(N1609), .B(N2989), .CI(N2457));
ADDFX1 inst_cellmath__43_0_I1188 (.CO(N3203), .S(N2775), .A(N2185), .B(N3302), .CI(N3031));
ADDFX1 inst_cellmath__43_0_I1189 (.CO(N2097), .S(N1669), .A(N2767), .B(N1916), .CI(N1652));
ADDFX1 inst_cellmath__43_0_I1190 (.CO(N2952), .S(N2529), .A(N3345), .B(N2500), .CI(N2229));
ADDFX1 inst_cellmath__43_0_I1191 (.CO(N1847), .S(N3380), .A(N1964), .B(N3073), .CI(N2813));
ADDFX1 inst_cellmath__43_0_I1192 (.CO(N2702), .S(N2272), .A(N2546), .B(N1700), .CI(N3393));
ADDFX1 inst_cellmath__43_0_I1193 (.CO(N1597), .S(N3130), .A(N2028), .B(N3140), .CI(N2887));
ADDFX1 inst_cellmath__43_0_I1194 (.CO(N2454), .S(N2019), .A(N2637), .B(N1780), .CI(N3491));
ADDFX1 inst_cellmath__43_0_I1195 (.CO(N3309), .S(N2878), .A(N3022), .B(N2389), .CI(N1918));
ADDFX1 inst_cellmath__43_0_I1196 (.CO(N2200), .S(N1771), .A(N1669), .B(N2775), .CI(N2529));
ADDFX1 inst_cellmath__43_0_I1197 (.CO(N3057), .S(N2628), .A(N2272), .B(N3380), .CI(N3243));
ADDFX1 inst_cellmath__43_0_I1198 (.CO(N1953), .S(N3482), .A(N2993), .B(N2136), .CI(N1884));
ADDFX1 inst_cellmath__43_0_I1199 (.CO(N2811), .S(N2382), .A(N3130), .B(N2742), .CI(N2019));
ADDFX1 inst_cellmath__43_0_I1200 (.CO(N1707), .S(N3234), .A(N2878), .B(N1639), .CI(N1771));
ADDFX1 inst_cellmath__43_0_I1201 (.CO(N2563), .S(N2127), .A(N2493), .B(N2628), .CI(N3348));
ADDFX1 inst_cellmath__43_0_I1202 (.CO(N3416), .S(N2985), .A(N2382), .B(N3482), .CI(N2242));
ADDFX1 inst_cellmath__43_0_I1203 (.CO(N2308), .S(N1877), .A(N3234), .B(N3093), .CI(N2127));
ADDFX1 inst_cellmath__43_0_I1204 (.CO(N3165), .S(N2735), .A(N2985), .B(N1990), .CI(N2849));
ADDFX1 inst_cellmath__43_0_I1205 (.CO(N2054), .S(N1630), .A(N1742), .B(N1877), .CI(N2735));
ADDFX1 inst_cellmath__43_0_I1206 (.CO(N2913), .S(N2485), .A(N1618), .B(N3381), .CI(N2465));
ADDFX1 inst_cellmath__43_0_I1207 (.CO(N1807), .S(N3340), .A(N3310), .B(N2730), .CI(N2193));
ADDFX1 inst_cellmath__43_0_I1208 (.CO(N2661), .S(N2233), .A(N1926), .B(N3041), .CI(N2774));
ADDFX1 inst_cellmath__43_0_I1209 (.CO(N1555), .S(N3086), .A(N2509), .B(N1662), .CI(N3354));
ADDFX1 inst_cellmath__43_0_I1210 (.CO(N2414), .S(N1983), .A(N3082), .B(N2236), .CI(N1973));
ADDFX1 inst_cellmath__43_0_I1211 (.CO(N3267), .S(N2840), .A(N1708), .B(N2819), .CI(N2555));
ADDFX1 inst_cellmath__43_0_I1212 (.CO(N2162), .S(N1736), .A(N2282), .B(N3403), .CI(N3453));
ADDFX1 inst_cellmath__43_0_I1213 (.CO(N3016), .S(N2591), .A(N3203), .B(N2348), .CI(N2097));
ADDFX1 inst_cellmath__43_0_I1214 (.CO(N1908), .S(N3446), .A(N1847), .B(N2952), .CI(N2702));
ADDFX1 inst_cellmath__43_0_I1215 (.CO(N2768), .S(N2340), .A(N3340), .B(N2485), .CI(N2233));
ADDFX1 inst_cellmath__43_0_I1216 (.CO(N1664), .S(N3195), .A(N1983), .B(N3086), .CI(N2840));
ADDFX1 inst_cellmath__43_0_I1217 (.CO(N2518), .S(N2087), .A(N2454), .B(N1597), .CI(N1736));
ADDFX1 inst_cellmath__43_0_I1218 (.CO(N3374), .S(N2944), .A(N2591), .B(N3309), .CI(N3446));
ADDFX1 inst_cellmath__43_0_I1219 (.CO(N2267), .S(N1838), .A(N3057), .B(N2200), .CI(N2340));
ADDFX1 inst_cellmath__43_0_I1220 (.CO(N3118), .S(N2695), .A(N1953), .B(N3195), .CI(N2811));
ADDFX1 inst_cellmath__43_0_I1221 (.CO(N2014), .S(N1590), .A(N2944), .B(N2087), .CI(N1707));
ADDFX1 inst_cellmath__43_0_I1222 (.CO(N2872), .S(N2445), .A(N1838), .B(N2563), .CI(N2695));
ADDFX1 inst_cellmath__43_0_I1223 (.CO(N1761), .S(N3300), .A(N1590), .B(N3416), .CI(N2308));
ADDFX1 inst_cellmath__43_0_I1224 (.CO(N2622), .S(N2192), .A(N3165), .B(N2445), .CI(N3300));
ADDFX1 inst_cellmath__43_0_I1225 (.CO(N3474), .S(N3046), .A(N3318), .B(N2273), .CI(N2205));
ADDFX1 inst_cellmath__43_0_I1226 (.CO(N2373), .S(N1944), .A(N3049), .B(N2474), .CI(N1936));
ADDFX1 inst_cellmath__43_0_I1227 (.CO(N3226), .S(N2800), .A(N1671), .B(N2784), .CI(N2519));
ADDFX1 inst_cellmath__43_0_I1228 (.CO(N2118), .S(N1698), .A(N2246), .B(N3364), .CI(N3092));
ADDFX1 inst_cellmath__43_0_I1229 (.CO(N2975), .S(N2553), .A(N2828), .B(N1981), .CI(N1715));
ADDFX1 inst_cellmath__43_0_I1230 (.CO(N1869), .S(N3407), .A(N3411), .B(N2565), .CI(N2291));
ADDFX1 inst_cellmath__43_0_I1231 (.CO(N2725), .S(N2298), .A(N2913), .B(N3138), .CI(N1807));
ADDFX1 inst_cellmath__43_0_I1232 (.CO(N1622), .S(N3155), .A(N1555), .B(N2661), .CI(N2414));
ADDFX1 inst_cellmath__43_0_I1233 (.CO(N2478), .S(N2042), .A(N3046), .B(N3267), .CI(N1944));
ADDFX1 inst_cellmath__43_0_I1234 (.CO(N3330), .S(N2903), .A(N1698), .B(N2800), .CI(N2553));
ADDFX1 inst_cellmath__43_0_I1235 (.CO(N2224), .S(N1796), .A(N2162), .B(N3407), .CI(N3016));
ADDFX1 inst_cellmath__43_0_I1236 (.CO(N3078), .S(N2653), .A(N2768), .B(N1908), .CI(N2298));
ADDFX1 inst_cellmath__43_0_I1237 (.CO(N1974), .S(N3510), .A(N3155), .B(N1664), .CI(N2042));
ADDFX1 inst_cellmath__43_0_I1238 (.CO(N2833), .S(N2404), .A(N2518), .B(N2903), .CI(N1796));
ADDFX1 inst_cellmath__43_0_I1239 (.CO(N1728), .S(N3257), .A(N2267), .B(N3374), .CI(N2653));
ADDFX1 inst_cellmath__43_0_I1240 (.CO(N2582), .S(N2153), .A(N3510), .B(N3118), .CI(N2404));
ADDFX1 inst_cellmath__43_0_I1241 (.CO(N3438), .S(N3007), .A(N3257), .B(N2014), .CI(N2872));
ADDFX1 inst_cellmath__43_0_I1242 (.CO(N2331), .S(N1898), .A(N1761), .B(N2153), .CI(N3007));
ADDFX1 inst_cellmath__43_0_I1243 (.CO(N3185), .S(N2760), .A(N3059), .B(N3127), .CI(N1947));
ADDFX1 inst_cellmath__43_0_I1244 (.CO(N2079), .S(N1654), .A(N2794), .B(N2211), .CI(N1681));
ADDFX1 inst_cellmath__43_0_I1245 (.CO(N2934), .S(N2507), .A(N3372), .B(N2527), .CI(N2255));
ADDFX1 inst_cellmath__43_0_I1246 (.CO(N1828), .S(N3366), .A(N1987), .B(N3101), .CI(N2838));
ADDFX1 inst_cellmath__43_0_I1247 (.CO(N2686), .S(N2257), .A(N2572), .B(N1723), .CI(N3419));
ADDFX1 inst_cellmath__43_0_I1248 (.CO(N1580), .S(N3109), .A(N3147), .B(N2300), .CI(N2029));
ADDFX1 inst_cellmath__43_0_I1249 (.CO(N2438), .S(N2007), .A(N2373), .B(N3474), .CI(N3226));
ADDFX1 inst_cellmath__43_0_I1250 (.CO(N3292), .S(N2863), .A(N2975), .B(N2118), .CI(N1869));
ADDFX1 inst_cellmath__43_0_I1251 (.CO(N2183), .S(N1753), .A(N1654), .B(N2760), .CI(N2507));
ADDFX1 inst_cellmath__43_0_I1252 (.CO(N3036), .S(N2615), .A(N2257), .B(N3366), .CI(N3109));
ADDFX1 inst_cellmath__43_0_I1253 (.CO(N1934), .S(N3468), .A(N1622), .B(N2725), .CI(N2478));
ADDFX1 inst_cellmath__43_0_I1254 (.CO(N2792), .S(N2363), .A(N2007), .B(N3330), .CI(N2863));
ADDFX1 inst_cellmath__43_0_I1255 (.CO(N1686), .S(N3219), .A(N1753), .B(N2224), .CI(N2615));
ADDFX1 inst_cellmath__43_0_I1256 (.CO(N2545), .S(N2111), .A(N1974), .B(N3078), .CI(N2363));
ADDFX1 inst_cellmath__43_0_I1257 (.CO(N3399), .S(N2965), .A(N2833), .B(N3468), .CI(N3219));
ADDFX1 inst_cellmath__43_0_I1258 (.CO(N2286), .S(N1862), .A(N2111), .B(N1728), .CI(N2582));
ADDFX1 inst_cellmath__43_0_I1259 (.CO(N3146), .S(N2716), .A(N3438), .B(N2965), .CI(N1862));
ADDFX1 inst_cellmath__43_0_I1260 (.CO(N2034), .S(N1611), .A(N2803), .B(N2020), .CI(N1692));
ADDFX1 inst_cellmath__43_0_I1261 (.CO(N2894), .S(N2469), .A(N2537), .B(N1954), .CI(N3379));
ADDFX1 inst_cellmath__43_0_I1262 (.CO(N1785), .S(N3323), .A(N3111), .B(N2265), .CI(N1997));
ADDFX1 inst_cellmath__43_0_I1263 (.CO(N2642), .S(N2215), .A(N1733), .B(N2844), .CI(N2581));
ADDFX1 inst_cellmath__43_0_I1264 (.CO(N3500), .S(N3069), .A(N2309), .B(N3425), .CI(N3159));
ADDFX1 inst_cellmath__43_0_I1265 (.CO(N2395), .S(N1965), .A(N2888), .B(N2038), .CI(N3185));
ADDFX1 inst_cellmath__43_0_I1266 (.CO(N3248), .S(N2823), .A(N2934), .B(N2079), .CI(N1828));
ADDFX1 inst_cellmath__43_0_I1267 (.CO(N2143), .S(N1719), .A(N1580), .B(N2686), .CI(N1611));
ADDFX1 inst_cellmath__43_0_I1268 (.CO(N2997), .S(N2574), .A(N3323), .B(N2469), .CI(N2215));
ADDFX1 inst_cellmath__43_0_I1269 (.CO(N1889), .S(N3429), .A(N2438), .B(N3069), .CI(N3292));
ADDFX1 inst_cellmath__43_0_I1270 (.CO(N2750), .S(N2322), .A(N2183), .B(N1965), .CI(N2823));
ADDFX1 inst_cellmath__43_0_I1271 (.CO(N1644), .S(N3175), .A(N1719), .B(N3036), .CI(N2574));
ADDFX1 inst_cellmath__43_0_I1272 (.CO(N2498), .S(N2069), .A(N2792), .B(N1934), .CI(N3429));
ADDFX1 inst_cellmath__43_0_I1273 (.CO(N3356), .S(N2924), .A(N1686), .B(N2322), .CI(N3175));
ADDFX1 inst_cellmath__43_0_I1274 (.CO(N2247), .S(N1818), .A(N2069), .B(N2545), .CI(N3399));
ADDFX1 inst_cellmath__43_0_I1275 (.CO(N3099), .S(N2677), .A(N2286), .B(N2924), .CI(N1818));
ADDFX1 inst_cellmath__43_0_I1276 (.CO(N1998), .S(N1569), .A(N2547), .B(N2879), .CI(N3391));
ADDFX1 inst_cellmath__43_0_I1277 (.CO(N2854), .S(N2428), .A(N2274), .B(N1701), .CI(N3119));
ADDFX1 inst_cellmath__43_0_I1278 (.CO(N1745), .S(N3282), .A(N2853), .B(N2005), .CI(N1741));
ADDFX1 inst_cellmath__43_0_I1279 (.CO(N2605), .S(N2174), .A(N3434), .B(N2590), .CI(N2318));
ADDFX1 inst_cellmath__43_0_I1280 (.CO(N3459), .S(N3028), .A(N2048), .B(N3167), .CI(N2896));
ADDFX1 inst_cellmath__43_0_I1281 (.CO(N2355), .S(N1924), .A(N2034), .B(N1779), .CI(N2894));
ADDFX1 inst_cellmath__43_0_I1282 (.CO(N3211), .S(N2782), .A(N2642), .B(N1785), .CI(N3500));
ADDFX1 inst_cellmath__43_0_I1283 (.CO(N2103), .S(N1676), .A(N2428), .B(N1569), .CI(N3282));
ADDFX1 inst_cellmath__43_0_I1284 (.CO(N2957), .S(N2535), .A(N3028), .B(N2174), .CI(N2395));
ADDFX1 inst_cellmath__43_0_I1285 (.CO(N1853), .S(N3389), .A(N2143), .B(N3248), .CI(N2997));
ADDFX1 inst_cellmath__43_0_I1286 (.CO(N2708), .S(N2279), .A(N2782), .B(N1924), .CI(N1889));
ADDFX1 inst_cellmath__43_0_I1287 (.CO(N1603), .S(N3137), .A(N2535), .B(N1676), .CI(N2750));
ADDFX1 inst_cellmath__43_0_I1288 (.CO(N2461), .S(N2026), .A(N1644), .B(N3389), .CI(N2279));
ADDFX1 inst_cellmath__43_0_I1289 (.CO(N3315), .S(N2885), .A(N3137), .B(N2498), .CI(N3356));
ADDFX1 inst_cellmath__43_0_I1290 (.CO(N2206), .S(N1778), .A(N2247), .B(N2026), .CI(N2885));
ADDFX1 inst_cellmath__43_0_I1291 (.CO(N3063), .S(N2635), .A(N2283), .B(N1769), .CI(N3128));
ADDFX1 inst_cellmath__43_0_I1292 (.CO(N1958), .S(N3487), .A(N2012), .B(N3401), .CI(N2861));
ADDFX1 inst_cellmath__43_0_I1293 (.CO(N2814), .S(N2387), .A(N2595), .B(N1747), .CI(N3442));
ADDFX1 inst_cellmath__43_0_I1294 (.CO(N1712), .S(N3241), .A(N3174), .B(N2326), .CI(N2057));
ADDFX1 inst_cellmath__43_0_I1295 (.CO(N2566), .S(N2131), .A(N1787), .B(N2904), .CI(N2638));
ADDFX1 inst_cellmath__43_0_I1296 (.CO(N3420), .S(N2990), .A(N2854), .B(N1998), .CI(N1745));
ADDFX1 inst_cellmath__43_0_I1297 (.CO(N2314), .S(N1880), .A(N3459), .B(N2605), .CI(N2635));
ADDFX1 inst_cellmath__43_0_I1298 (.CO(N3168), .S(N2738), .A(N2387), .B(N3487), .CI(N3241));
ADDFX1 inst_cellmath__43_0_I1299 (.CO(N2060), .S(N1636), .A(N2355), .B(N2131), .CI(N3211));
ADDFX1 inst_cellmath__43_0_I1300 (.CO(N2916), .S(N2490), .A(N2990), .B(N2103), .CI(N2957));
ADDFX1 inst_cellmath__43_0_I1301 (.CO(N1810), .S(N3346), .A(N2738), .B(N1880), .CI(N1853));
ADDFX1 inst_cellmath__43_0_I1302 (.CO(N2667), .S(N2238), .A(N2708), .B(N1636), .CI(N2490));
ADDFX1 inst_cellmath__43_0_I1303 (.CO(N1559), .S(N3090), .A(N3346), .B(N1603), .CI(N2461));
ADDFX1 inst_cellmath__43_0_I1304 (.CO(N2418), .S(N1989), .A(N3315), .B(N2238), .CI(N3090));
ADDFX1 inst_cellmath__43_0_I1305 (.CO(N3273), .S(N2846), .A(N2018), .B(N2629), .CI(N2873));
ADDFX1 inst_cellmath__43_0_I1306 (.CO(N2166), .S(N1739), .A(N1755), .B(N3139), .CI(N2604));
ADDFX1 inst_cellmath__43_0_I1307 (.CO(N3020), .S(N2597), .A(N2338), .B(N3449), .CI(N3183));
ADDFX1 inst_cellmath__43_0_I1308 (.CO(N1914), .S(N3450), .A(N2914), .B(N2065), .CI(N1801));
ADDFX1 inst_cellmath__43_0_I1309 (.CO(N2772), .S(N2343), .A(N3492), .B(N2648), .CI(N3063));
ADDFX1 inst_cellmath__43_0_I1310 (.CO(N1667), .S(N3200), .A(N2814), .B(N1958), .CI(N1712));
ADDFX1 inst_cellmath__43_0_I1311 (.CO(N2525), .S(N2094), .A(N2846), .B(N2566), .CI(N1739));
ADDFX1 inst_cellmath__43_0_I1312 (.CO(N3377), .S(N2947), .A(N3450), .B(N2597), .CI(N3420));
ADDFX1 inst_cellmath__43_0_I1313 (.CO(N2270), .S(N1844), .A(N2314), .B(N2343), .CI(N3168));
ADDFX1 inst_cellmath__43_0_I1314 (.CO(N3126), .S(N2699), .A(N2094), .B(N3200), .CI(N2060));
ADDFX1 inst_cellmath__43_0_I1315 (.CO(N2016), .S(N1593), .A(N2916), .B(N2947), .CI(N1844));
ADDFX1 inst_cellmath__43_0_I1316 (.CO(N2876), .S(N2451), .A(N2699), .B(N1810), .CI(N2667));
ADDFX1 inst_cellmath__43_0_I1317 (.CO(N1768), .S(N3306), .A(N1559), .B(N1593), .CI(N2451));
ADDFX1 inst_cellmath__43_0_I1318 (.CO(N2626), .S(N2197), .A(N1762), .B(N3483), .CI(N2613));
ADDFX1 inst_cellmath__43_0_I1319 (.CO(N3479), .S(N3054), .A(N3457), .B(N2880), .CI(N2345));
ADDFX1 inst_cellmath__43_0_I1320 (.CO(N2379), .S(N1950), .A(N2074), .B(N3192), .CI(N2920));
ADDFX1 inst_cellmath__43_0_I1321 (.CO(N3232), .S(N2807), .A(N2658), .B(N1809), .CI(N3502));
ADDFX1 inst_cellmath__43_0_I1322 (.CO(N2124), .S(N1704), .A(N3273), .B(N2388), .CI(N2166));
ADDFX1 inst_cellmath__43_0_I1323 (.CO(N2982), .S(N2559), .A(N1914), .B(N3020), .CI(N2197));
ADDFX1 inst_cellmath__43_0_I1324 (.CO(N1875), .S(N3413), .A(N1950), .B(N3054), .CI(N2807));
ADDFX1 inst_cellmath__43_0_I1325 (.CO(N2731), .S(N2304), .A(N1667), .B(N2772), .CI(N2525));
ADDFX1 inst_cellmath__43_0_I1326 (.CO(N1627), .S(N3161), .A(N3377), .B(N1704), .CI(N2559));
ADDFX1 inst_cellmath__43_0_I1327 (.CO(N2483), .S(N2051), .A(N2270), .B(N3413), .CI(N2304));
ADDFX1 inst_cellmath__43_0_I1328 (.CO(N3336), .S(N2909), .A(N3161), .B(N3126), .CI(N2016));
ADDFX1 inst_cellmath__43_0_I1329 (.CO(N2230), .S(N1803), .A(N2876), .B(N2051), .CI(N2909));
ADDFX1 inst_cellmath__43_0_I1330 (.CO(N3083), .S(N2659), .A(N3466), .B(N2380), .CI(N2357));
ADDFX1 inst_cellmath__43_0_I1331 (.CO(N1979), .S(N1553), .A(N3199), .B(N2620), .CI(N2083));
ADDFX1 inst_cellmath__43_0_I1332 (.CO(N2839), .S(N2411), .A(N1816), .B(N2928), .CI(N2664));
ADDFX1 inst_cellmath__43_0_I1333 (.CO(N1734), .S(N3264), .A(N2397), .B(N3511), .CI(N3244));
ADDFX1 inst_cellmath__43_0_I1334 (.CO(N2588), .S(N2160), .A(N3479), .B(N2626), .CI(N2379));
ADDFX1 inst_cellmath__43_0_I1335 (.CO(N3443), .S(N3013), .A(N2659), .B(N3232), .CI(N1553));
ADDFX1 inst_cellmath__43_0_I1336 (.CO(N2336), .S(N1905), .A(N3264), .B(N2411), .CI(N2124));
ADDFX1 inst_cellmath__43_0_I1337 (.CO(N3193), .S(N2765), .A(N1875), .B(N2982), .CI(N2160));
ADDFX1 inst_cellmath__43_0_I1338 (.CO(N2084), .S(N1660), .A(N2731), .B(N3013), .CI(N1905));
ADDFX1 inst_cellmath__43_0_I1339 (.CO(N2939), .S(N2517), .A(N2765), .B(N1627), .CI(N2483));
ADDFX1 inst_cellmath__43_0_I1340 (.CO(N1836), .S(N3370), .A(N3336), .B(N1660), .CI(N2517));
ADDFX1 inst_cellmath__43_0_I1341 (.CO(N2691), .S(N2263), .A(N3209), .B(N3235), .CI(N2092));
ADDFX1 inst_cellmath__43_0_I1342 (.CO(N1585), .S(N3117), .A(N2941), .B(N2365), .CI(N1826));
ADDFX1 inst_cellmath__43_0_I1343 (.CO(N2444), .S(N2010), .A(N1556), .B(N2672), .CI(N2407));
ADDFX1 inst_cellmath__43_0_I1344 (.CO(N3296), .S(N2868), .A(N2137), .B(N3253), .CI(N3083));
ADDFX1 inst_cellmath__43_0_I1345 (.CO(N2188), .S(N1760), .A(N2839), .B(N1979), .CI(N1734));
ADDFX1 inst_cellmath__43_0_I1346 (.CO(N3043), .S(N2618), .A(N3117), .B(N2263), .CI(N2010));
ADDFX1 inst_cellmath__43_0_I1347 (.CO(N1939), .S(N3472), .A(N2868), .B(N2588), .CI(N3443));
ADDFX1 inst_cellmath__43_0_I1348 (.CO(N2797), .S(N2370), .A(N2336), .B(N1760), .CI(N2618));
ADDFX1 inst_cellmath__43_0_I1349 (.CO(N1694), .S(N3223), .A(N3472), .B(N3193), .CI(N2084));
ADDFX1 inst_cellmath__43_0_I1350 (.CO(N2549), .S(N2115), .A(N2939), .B(N2370), .CI(N3223));
ADDFX1 inst_cellmath__43_0_I1351 (.CO(N3404), .S(N2972), .A(N2949), .B(N2128), .CI(N1835));
ADDFX1 inst_cellmath__43_0_I1352 (.CO(N2293), .S(N1866), .A(N2681), .B(N2102), .CI(N1564));
ADDFX1 inst_cellmath__43_0_I1353 (.CO(N3150), .S(N2722), .A(N3262), .B(N2416), .CI(N2145));
ADDFX1 inst_cellmath__43_0_I1354 (.CO(N2039), .S(N1619), .A(N2691), .B(N2991), .CI(N1585));
ADDFX1 inst_cellmath__43_0_I1355 (.CO(N2898), .S(N2475), .A(N2972), .B(N2444), .CI(N1866));
ADDFX1 inst_cellmath__43_0_I1356 (.CO(N1791), .S(N3327), .A(N3296), .B(N2722), .CI(N2188));
ADDFX1 inst_cellmath__43_0_I1357 (.CO(N2650), .S(N2221), .A(N1619), .B(N3043), .CI(N2475));
ADDFX1 inst_cellmath__43_0_I1358 (.CO(N3505), .S(N3075), .A(N3327), .B(N1939), .CI(N2797));
ADDFX1 inst_cellmath__43_0_I1359 (.CO(N2400), .S(N1971), .A(N1694), .B(N2221), .CI(N3075));
ADDFX1 inst_cellmath__43_0_I1360 (.CO(N3255), .S(N2829), .A(N2690), .B(N2983), .CI(N1574));
ADDFX1 inst_cellmath__43_0_I1361 (.CO(N2149), .S(N1725), .A(N2426), .B(N1843), .CI(N3270));
ADDFX1 inst_cellmath__43_0_I1362 (.CO(N3003), .S(N2579), .A(N2999), .B(N2154), .CI(N1885));
ADDFX1 inst_cellmath__43_0_I1363 (.CO(N1896), .S(N3435), .A(N2293), .B(N3404), .CI(N3150));
ADDFX1 inst_cellmath__43_0_I1364 (.CO(N2756), .S(N2328), .A(N1725), .B(N2829), .CI(N2579));
ADDFX1 inst_cellmath__43_0_I1365 (.CO(N1650), .S(N3181), .A(N2898), .B(N2039), .CI(N3435));
ADDFX1 inst_cellmath__43_0_I1366 (.CO(N2505), .S(N2075), .A(N2328), .B(N1791), .CI(N2650));
ADDFX1 inst_cellmath__43_0_I1367 (.CO(N3362), .S(N2930), .A(N3505), .B(N3181), .CI(N2075));
ADDFX1 inst_cellmath__43_0_I1368 (.CO(N2253), .S(N1824), .A(N2436), .B(N1878), .CI(N3277));
ADDFX1 inst_cellmath__43_0_I1369 (.CO(N3107), .S(N2683), .A(N2163), .B(N1587), .CI(N3010));
ADDFX1 inst_cellmath__43_0_I1370 (.CO(N2003), .S(N1576), .A(N2743), .B(N1893), .CI(N3255));
ADDFX1 inst_cellmath__43_0_I1371 (.CO(N2859), .S(N2434), .A(N3003), .B(N2149), .CI(N1824));
ADDFX1 inst_cellmath__43_0_I1372 (.CO(N1750), .S(N3288), .A(N1896), .B(N2683), .CI(N1576));
ADDFX1 inst_cellmath__43_0_I1373 (.CO(N2610), .S(N2179), .A(N2434), .B(N2756), .CI(N1650));
ADDFX1 inst_cellmath__43_0_I1374 (.CO(N3464), .S(N3033), .A(N2505), .B(N3288), .CI(N2179));
ADDFX1 inst_cellmath__43_0_I1375 (.CO(N2362), .S(N1929), .A(N2170), .B(N2736), .CI(N3018));
ADDFX1 inst_cellmath__43_0_I1376 (.CO(N3215), .S(N2788), .A(N1903), .B(N3286), .CI(N2751));
ADDFX1 inst_cellmath__43_0_I1377 (.CO(N2108), .S(N1684), .A(N2253), .B(N1638), .CI(N3107));
ADDFX1 inst_cellmath__43_0_I1378 (.CO(N2964), .S(N2540), .A(N2788), .B(N1929), .CI(N2003));
ADDFX1 inst_cellmath__43_0_I1379 (.CO(N1858), .S(N3395), .A(N1684), .B(N2859), .CI(N1750));
ADDFX1 inst_cellmath__43_0_I1380 (.CO(N2712), .S(N2285), .A(N2610), .B(N2540), .CI(N3395));
ADDFX1 inst_cellmath__43_0_I1381 (.CO(N1610), .S(N3141), .A(N1911), .B(N1628), .CI(N2761));
ADDFX1 inst_cellmath__43_0_I1382 (.CO(N2466), .S(N2030), .A(N1647), .B(N3026), .CI(N2494));
ADDFX1 inst_cellmath__43_0_I1383 (.CO(N3319), .S(N2890), .A(N3215), .B(N2362), .CI(N3141));
ADDFX1 inst_cellmath__43_0_I1384 (.CO(N2212), .S(N1781), .A(N2108), .B(N2030), .CI(N2964));
ADDFX1 inst_cellmath__43_0_I1385 (.CO(N3066), .S(N2639), .A(N1858), .B(N2890), .CI(N1781));
ADDFX1 inst_cellmath__43_0_I1386 (.CO(N1962), .S(N3495), .A(N1657), .B(N2486), .CI(N2502));
ADDFX1 inst_cellmath__43_0_I1387 (.CO(N2820), .S(N2390), .A(N3349), .B(N2769), .CI(N1610));
ADDFX1 inst_cellmath__43_0_I1388 (.CO(N1716), .S(N3245), .A(N3495), .B(N2466), .CI(N2390));
ADDFX1 inst_cellmath__43_0_I1389 (.CO(N2570), .S(N2139), .A(N2212), .B(N3319), .CI(N3245));
ADDFX1 inst_cellmath__43_0_I1390 (.CO(N3426), .S(N2994), .A(N3357), .B(N3341), .CI(N2240));
ADDFX1 inst_cellmath__43_0_I1391 (.CO(N2319), .S(N1887), .A(N1962), .B(N2512), .CI(N2994));
ADDFX1 inst_cellmath__43_0_I1392 (.CO(N3172), .S(N2746), .A(N1887), .B(N2820), .CI(N1716));
ADDFX1 inst_cellmath__43_0_I1393 (.CO(N2066), .S(N1641), .A(N3094), .B(N2231), .CI(N2250));
ADDFX1 inst_cellmath__43_0_I1394 (.CO(N2921), .S(N2496), .A(N1641), .B(N3426), .CI(N2319));
ADDFX1 inst_cellmath__43_0_I1395 (.CO(N2159), .S(N3352), .A(N1991), .B(N3087), .CI(N2066));
OR4X1 inst_cellmath__43_0_I9658 (.Y(N2244), .A(N3303), .B(N1798), .C(N3335), .D(N1765));
NOR2XL inst_cellmath__43_0_I1397 (.Y(N2673), .A(N3184), .B(N1945));
NAND2XL inst_cellmath__43_0_I1398 (.Y(N3097), .A(N3184), .B(N1945));
AND2XL inst_cellmath__43_0_I1400 (.Y(N1995), .A(N2801), .B(N1695));
NOR2XL inst_cellmath__43_0_I1401 (.Y(N2424), .A(N3408), .B(N2294));
NAND2XL inst_cellmath__43_0_I1402 (.Y(N2851), .A(N3408), .B(N2294));
AND2XL inst_cellmath__43_0_I1404 (.Y(N1584), .A(N2726), .B(N1797));
NOR2XL inst_cellmath__43_0_I1405 (.Y(N2171), .A(N2222), .B(N2150));
NAND2XL inst_cellmath__43_0_I1406 (.Y(N2602), .A(N2222), .B(N2150));
AND2XL inst_cellmath__43_0_I1408 (.Y(N3455), .A(N2583), .B(N3363));
NOR2XL inst_cellmath__43_0_I1409 (.Y(N1920), .A(N1829), .B(N3469));
NAND2XL inst_cellmath__43_0_I1410 (.Y(N2352), .A(N1829), .B(N3469));
NOR2XL inst_cellmath__43_0_I1411 (.Y(N2778), .A(N1931), .B(N2470));
NOR2XL inst_cellmath__43_0_I1413 (.Y(N1673), .A(N2891), .B(N2323));
NAND2XL inst_cellmath__43_0_I1414 (.Y(N2100), .A(N2891), .B(N2323));
NOR2XL inst_cellmath__43_0_I1415 (.Y(N2532), .A(N2747), .B(N3029));
NAND2XL inst_cellmath__43_0_I1416 (.Y(N2955), .A(N2747), .B(N3029));
NOR2XL inst_cellmath__43_0_I1417 (.Y(N3384), .A(N3460), .B(N2636));
NAND2XL inst_cellmath__43_0_I1418 (.Y(N1851), .A(N3460), .B(N2636));
NOR2XL inst_cellmath__43_0_I1419 (.Y(N2276), .A(N3062), .B(N3091));
NOR2XL inst_cellmath__43_0_I1421 (.Y(N3133), .A(N1560), .B(N2450));
NAND2XL inst_cellmath__43_0_I1422 (.Y(N1599), .A(N1560), .B(N2450));
NOR2XL inst_cellmath__43_0_I1423 (.Y(N2022), .A(N2877), .B(N2660));
NAND2XL inst_cellmath__43_0_I1424 (.Y(N2459), .A(N2877), .B(N2660));
NOR2XL inst_cellmath__43_0_I1425 (.Y(N2882), .A(N3084), .B(N1758));
NAND2XL inst_cellmath__43_0_I1426 (.Y(N3312), .A(N3084), .B(N1758));
AOI21XL inst_cellmath__43_0_I1427 (.Y(N2631), .A0(N3097), .A1(N2244), .B0(N2673));
OAI22XL inst_cellmath__43_0_I3427 (.Y(N2130), .A0(N1995), .A1(N2631), .B0(N2801), .B1(N1695));
AOI21XL inst_cellmath__43_0_I1431 (.Y(N1632), .A0(N2851), .A1(N2130), .B0(N2424));
OAI22XL inst_cellmath__43_0_I3428 (.Y(N2842), .A0(N1584), .A1(N1632), .B0(N2726), .B1(N1797));
AOI21XL inst_cellmath__43_0_I1434 (.Y(N2090), .A0(N2602), .A1(N2842), .B0(N2171));
OAI22XL inst_cellmath__43_0_I3429 (.Y(N3051), .A0(N3455), .A1(N2090), .B0(N2583), .B1(N3363));
AOI21XL inst_cellmath__43_0_I1438 (.Y(N2046), .A0(N2352), .A1(N3051), .B0(N1920));
AOI21XL inst_cellmath__43_0_I1439 (.Y(N1799), .A0(N2100), .A1(N2778), .B0(N1673));
OAI2BB1X1 inst_cellmath__43_0_I3430 (.Y(N2226), .A0N(N1931), .A1N(N2470), .B0(N2100));
OAI21XL inst_cellmath__43_0_I1441 (.Y(N2514), .A0(N2226), .A1(N2046), .B0(N1799));
AOI21XL inst_cellmath__43_0_I1442 (.Y(N2259), .A0(N1851), .A1(N2532), .B0(N3384));
INVXL inst_cellmath__43_0_I1443 (.Y(N3104), .A(N2259));
AOI31X1 inst_cellmath__43_0_I1445 (.Y(N2471), .A0(N1851), .A1(N2955), .A2(N2514), .B0(N3104));
AOI21XL inst_cellmath__43_0_I1446 (.Y(N2217), .A0(N1599), .A1(N2276), .B0(N3133));
OAI2BB1X1 inst_cellmath__43_0_I3431 (.Y(N2646), .A0N(N3062), .A1N(N3091), .B0(N1599));
OAI21XL inst_cellmath__43_0_I1448 (.Y(N2432), .A0(N2646), .A1(N2471), .B0(N2217));
AO21XL inst_cellmath__43_0_I1449 (.Y(N1961), .A0(N3312), .A1(N2022), .B0(N2882));
AOI31X1 inst_cellmath__43_0_I1455 (.Y(N1883), .A0(N3312), .A1(N2459), .A2(N2432), .B0(N1961));
NOR2XL inst_cellmath__43_0_I1490 (.Y(N3373), .A(N2147), .B(N2541));
XOR2XL inst_cellmath__43_0_I1491 (.Y(N1839), .A(N2147), .B(N2541));
NOR2XL inst_cellmath__43_0_I1492 (.Y(N2266), .A(N2961), .B(N2245));
XOR2XL inst_cellmath__43_0_I1493 (.Y(N2694), .A(N2961), .B(N2245));
NOR2XL inst_cellmath__43_0_I1494 (.Y(N3120), .A(N2671), .B(N2812));
XOR2XL inst_cellmath__43_0_I1495 (.Y(N1589), .A(N2671), .B(N2812));
NOR2XL inst_cellmath__43_0_I1496 (.Y(N2013), .A(N3237), .B(N2268));
XOR2XL inst_cellmath__43_0_I1497 (.Y(N2447), .A(N3237), .B(N2268));
NOR2XL inst_cellmath__43_0_I1498 (.Y(N2871), .A(N2697), .B(N3441));
XOR2XL inst_cellmath__43_0_I1499 (.Y(N3299), .A(N2697), .B(N3441));
NOR2XL inst_cellmath__43_0_I1500 (.Y(N1763), .A(N1902), .B(N2647));
XOR2XL inst_cellmath__43_0_I1501 (.Y(N2191), .A(N1902), .B(N2647));
NOR2XL inst_cellmath__43_0_I1502 (.Y(N2621), .A(N3072), .B(N1854));
XOR2XL inst_cellmath__43_0_I1503 (.Y(N3045), .A(N3072), .B(N1854));
NOR2XL inst_cellmath__43_0_I1504 (.Y(N3475), .A(N2281), .B(N2169));
XOR2XL inst_cellmath__43_0_I1505 (.Y(N1943), .A(N2281), .B(N2169));
NOR2XL inst_cellmath__43_0_I1506 (.Y(N2372), .A(N2598), .B(N1630));
XOR2XL inst_cellmath__43_0_I1507 (.Y(N2802), .A(N2598), .B(N1630));
NOR2XL inst_cellmath__43_0_I1508 (.Y(N3225), .A(N2054), .B(N2192));
XOR2XL inst_cellmath__43_0_I1509 (.Y(N1697), .A(N2054), .B(N2192));
NOR2XL inst_cellmath__43_0_I1510 (.Y(N2120), .A(N2622), .B(N1898));
XOR2XL inst_cellmath__43_0_I1511 (.Y(N2552), .A(N2622), .B(N1898));
NOR2XL inst_cellmath__43_0_I1512 (.Y(N2974), .A(N2331), .B(N2716));
XOR2XL inst_cellmath__43_0_I1513 (.Y(N3409), .A(N2331), .B(N2716));
NOR2XL inst_cellmath__43_0_I1514 (.Y(N1868), .A(N3146), .B(N2677));
XOR2XL inst_cellmath__43_0_I1515 (.Y(N2297), .A(N3146), .B(N2677));
NOR2XL inst_cellmath__43_0_I1516 (.Y(N2727), .A(N3099), .B(N1778));
XOR2XL inst_cellmath__43_0_I1517 (.Y(N3154), .A(N3099), .B(N1778));
NOR2XL inst_cellmath__43_0_I1518 (.Y(N1621), .A(N2206), .B(N1989));
XOR2XL inst_cellmath__43_0_I1519 (.Y(N2045), .A(N2206), .B(N1989));
NOR2XL inst_cellmath__43_0_I1520 (.Y(N2477), .A(N2418), .B(N3306));
XOR2XL inst_cellmath__43_0_I1521 (.Y(N2902), .A(N2418), .B(N3306));
NOR2XL inst_cellmath__43_0_I1522 (.Y(N3332), .A(N1768), .B(N1803));
XOR2XL inst_cellmath__43_0_I1523 (.Y(N1795), .A(N1768), .B(N1803));
NOR2XL inst_cellmath__43_0_I1524 (.Y(N2223), .A(N2230), .B(N3370));
XOR2XL inst_cellmath__43_0_I1525 (.Y(N2656), .A(N2230), .B(N3370));
NOR2XL inst_cellmath__43_0_I1526 (.Y(N3077), .A(N1836), .B(N2115));
XOR2XL inst_cellmath__43_0_I1527 (.Y(N3509), .A(N1836), .B(N2115));
NOR2XL inst_cellmath__43_0_I1528 (.Y(N1976), .A(N2549), .B(N1971));
XOR2XL inst_cellmath__43_0_I1529 (.Y(N2403), .A(N2549), .B(N1971));
NOR2XL inst_cellmath__43_0_I1530 (.Y(N2832), .A(N2400), .B(N2930));
XOR2XL inst_cellmath__43_0_I1531 (.Y(N3260), .A(N2400), .B(N2930));
NOR2XL inst_cellmath__43_0_I1532 (.Y(N1727), .A(N3362), .B(N3033));
XOR2XL inst_cellmath__43_0_I1533 (.Y(N2152), .A(N3362), .B(N3033));
NOR2XL inst_cellmath__43_0_I1534 (.Y(N2584), .A(N3464), .B(N2285));
XOR2XL inst_cellmath__43_0_I1535 (.Y(N3006), .A(N3464), .B(N2285));
NOR2XL inst_cellmath__43_0_I1536 (.Y(N3437), .A(N2712), .B(N2639));
XOR2XL inst_cellmath__43_0_I1537 (.Y(N1901), .A(N2712), .B(N2639));
NOR2XL inst_cellmath__43_0_I1538 (.Y(N2330), .A(N3066), .B(N2139));
XOR2XL inst_cellmath__43_0_I1539 (.Y(N2759), .A(N3066), .B(N2139));
NOR2XL inst_cellmath__43_0_I1540 (.Y(N3187), .A(N2746), .B(N2570));
XOR2XL inst_cellmath__43_0_I1541 (.Y(N1653), .A(N2746), .B(N2570));
NOR2XL inst_cellmath__43_0_I1542 (.Y(N2078), .A(N2496), .B(N3172));
XOR2XL inst_cellmath__43_0_I1543 (.Y(N2510), .A(N2496), .B(N3172));
NOR2XL inst_cellmath__43_0_I1544 (.Y(N2933), .A(N3352), .B(N2921));
XOR2XL inst_cellmath__43_0_I1545 (.Y(N3365), .A(N3352), .B(N2921));
OR2XL cmp_A_I9661 (.Y(N16704), .A(N2189), .B(N1726));
AO22XL cmp_A_I9662 (.Y(N2256), .A0(N16704), .A1(N1883), .B0(N2189), .B1(N1726));
AOI21XL inst_cellmath__43_0_I1547 (.Y(N3112), .A0(N2694), .A1(N3373), .B0(N2266));
NAND2XL inst_cellmath__43_0_I1548 (.Y(N1579), .A(N2694), .B(N1839));
AOI21XL inst_cellmath__43_0_I1549 (.Y(N2006), .A0(N2447), .A1(N3120), .B0(N2013));
NAND2XL inst_cellmath__43_0_I1550 (.Y(N2440), .A(N2447), .B(N1589));
AOI21XL inst_cellmath__43_0_I1551 (.Y(N2862), .A0(N2191), .A1(N2871), .B0(N1763));
NAND2XL inst_cellmath__43_0_I1552 (.Y(N3291), .A(N2191), .B(N3299));
AOI21XL inst_cellmath__43_0_I1553 (.Y(N1756), .A0(N1943), .A1(N2621), .B0(N3475));
NAND2XL inst_cellmath__43_0_I1554 (.Y(N2182), .A(N1943), .B(N3045));
AOI21XL inst_cellmath__43_0_I1555 (.Y(N2614), .A0(N1697), .A1(N2372), .B0(N3225));
NAND2XL inst_cellmath__43_0_I1556 (.Y(N3038), .A(N1697), .B(N2802));
AOI21XL inst_cellmath__43_0_I1557 (.Y(N3467), .A0(N3409), .A1(N2120), .B0(N2974));
NAND2XL inst_cellmath__43_0_I1558 (.Y(N1933), .A(N3409), .B(N2552));
AOI21XL inst_cellmath__43_0_I1559 (.Y(N2366), .A0(N3154), .A1(N1868), .B0(N2727));
NAND2XL inst_cellmath__43_0_I1560 (.Y(N2791), .A(N3154), .B(N2297));
AOI21XL inst_cellmath__43_0_I1561 (.Y(N3218), .A0(N2902), .A1(N1621), .B0(N2477));
NAND2XL inst_cellmath__43_0_I1562 (.Y(N1689), .A(N2902), .B(N2045));
AOI21XL inst_cellmath__43_0_I1563 (.Y(N2110), .A0(N2656), .A1(N3332), .B0(N2223));
NAND2XL inst_cellmath__43_0_I1564 (.Y(N2544), .A(N2656), .B(N1795));
AOI21XL inst_cellmath__43_0_I1565 (.Y(N2967), .A0(N2403), .A1(N3077), .B0(N1976));
NAND2XL inst_cellmath__43_0_I1566 (.Y(N3398), .A(N2403), .B(N3509));
AOI21XL inst_cellmath__43_0_I1567 (.Y(N1861), .A0(N2152), .A1(N2832), .B0(N1727));
NAND2XL inst_cellmath__43_0_I1568 (.Y(N2289), .A(N2152), .B(N3260));
AOI21XL inst_cellmath__43_0_I1569 (.Y(N2715), .A0(N1901), .A1(N2584), .B0(N3437));
NAND2XL inst_cellmath__43_0_I1570 (.Y(N3145), .A(N1901), .B(N3006));
AOI21XL inst_cellmath__43_0_I1571 (.Y(N1613), .A0(N1653), .A1(N2330), .B0(N3187));
NAND2XL inst_cellmath__43_0_I1572 (.Y(N2033), .A(N1653), .B(N2759));
AOI21XL inst_cellmath__43_0_I1573 (.Y(N2468), .A0(N3365), .A1(N2078), .B0(N2933));
OAI21XL inst_cellmath__43_0_I1574 (.Y(N3322), .A0(N1579), .A1(N2256), .B0(N3112));
OAI21XL inst_cellmath__43_0_I1575 (.Y(N2214), .A0(N3291), .A1(N2006), .B0(N2862));
NOR2XL inst_cellmath__43_0_I1576 (.Y(N2645), .A(N3291), .B(N2440));
OAI21XL inst_cellmath__43_0_I1577 (.Y(N3068), .A0(N3038), .A1(N1756), .B0(N2614));
NOR2XL inst_cellmath__43_0_I1578 (.Y(N3499), .A(N3038), .B(N2182));
OAI21XL inst_cellmath__43_0_I1579 (.Y(N1967), .A0(N2791), .A1(N3467), .B0(N2366));
NOR2XL inst_cellmath__43_0_I1580 (.Y(N2394), .A(N2791), .B(N1933));
OAI21XL inst_cellmath__43_0_I1581 (.Y(N2822), .A0(N2544), .A1(N3218), .B0(N2110));
NOR2XL inst_cellmath__43_0_I1582 (.Y(N3251), .A(N2544), .B(N1689));
OAI21XL inst_cellmath__43_0_I1583 (.Y(N1718), .A0(N2289), .A1(N2967), .B0(N1861));
NOR2XL inst_cellmath__43_0_I1584 (.Y(N2142), .A(N2289), .B(N3398));
AOI21XL inst_cellmath__43_0_I1585 (.Y(N3428), .A0(N2645), .A1(N3322), .B0(N2214));
AOI21XL inst_cellmath__43_0_I1586 (.Y(N2321), .A0(N2394), .A1(N3068), .B0(N1967));
NAND2XL inst_cellmath__43_0_I1587 (.Y(N2749), .A(N2394), .B(N3499));
AOI21XL inst_cellmath__43_0_I1588 (.Y(N3177), .A0(N2142), .A1(N2822), .B0(N1718));
OAI21XL inst_cellmath__43_0_I1589 (.Y(N2068), .A0(N2749), .A1(N3428), .B0(N2321));
INVXL inst_cellmath__43_0_I1590 (.Y(N3355), .A(N3177));
AOI31X1 inst_cellmath__43_0_I1591 (.Y(N1820), .A0(N2142), .A1(N3251), .A2(N2068), .B0(N3355));
INVXL inst_cellmath__43_0_I1592 (.Y(N2676), .A(N3499));
INVXL inst_cellmath__43_0_I1593 (.Y(N3102), .A(N3068));
OAI21XL inst_cellmath__43_0_I1594 (.Y(N1568), .A0(N2676), .A1(N3428), .B0(N3102));
INVXL inst_cellmath__43_0_I1595 (.Y(N1814), .A(N2068));
AOI21XL inst_cellmath__43_0_I1596 (.Y(N3281), .A0(N3251), .A1(N2068), .B0(N2822));
INVXL inst_cellmath__43_0_I1597 (.Y(N2241), .A(N1820));
OA21X1 inst_cellmath__43_0_I1598 (.Y(N3458), .A0(N2033), .A1(N2715), .B0(N1613));
OAI31X1 inst_cellmath__43_0_I1599 (.Y(N1923), .A0(N2033), .A1(N3145), .A2(N1820), .B0(N3458));
INVXL inst_cellmath__43_0_I1600 (.Y(N2781), .A(N2440));
INVXL inst_cellmath__43_0_I1601 (.Y(N3210), .A(N2006));
AOI21XL inst_cellmath__43_0_I1602 (.Y(N1678), .A0(N2781), .A1(N3322), .B0(N3210));
INVXL inst_cellmath__43_0_I1603 (.Y(N2670), .A(N3428));
OAI21XL inst_cellmath__43_0_I1604 (.Y(N3388), .A0(N2182), .A1(N3428), .B0(N1756));
INVXL inst_cellmath__43_0_I1605 (.Y(N3095), .A(N1568));
INVXL inst_cellmath__43_0_I1606 (.Y(N3136), .A(N1933));
INVXL inst_cellmath__43_0_I1607 (.Y(N1605), .A(N3467));
AOI21XL inst_cellmath__43_0_I1608 (.Y(N2025), .A0(N3136), .A1(N1568), .B0(N1605));
INVXL inst_cellmath__43_0_I1609 (.Y(N1562), .A(N1814));
OAI21XL inst_cellmath__43_0_I1610 (.Y(N1777), .A0(N1689), .A1(N1814), .B0(N3218));
INVXL inst_cellmath__43_0_I1611 (.Y(N1992), .A(N3281));
OAI21XL inst_cellmath__43_0_I1612 (.Y(N3490), .A0(N3398), .A1(N3281), .B0(N2967));
INVXL inst_cellmath__43_0_I1613 (.Y(N2423), .A(N2241));
INVXL inst_cellmath__43_0_I1614 (.Y(N3240), .A(N3145));
INVXL inst_cellmath__43_0_I1615 (.Y(N1711), .A(N2715));
AOI21XL inst_cellmath__43_0_I1616 (.Y(N2135), .A0(N3240), .A1(N2241), .B0(N1711));
INVXL inst_cellmath__43_0_I1617 (.Y(N2848), .A(N1923));
INVXL inst_cellmath__43_0_I1618 (.Y(N2313), .A(N2468));
AOI31X1 inst_cellmath__43_0_I1619 (.Y(N2741), .A0(N3365), .A1(N2510), .A2(N1923), .B0(N2313));
INVXL inst_cellmath__43_0_I1624 (.Y(N1988), .A(N3299));
INVXL inst_cellmath__43_0_I1625 (.Y(N2420), .A(N2871));
OAI21XL inst_cellmath__43_0_I1626 (.Y(N2845), .A0(N1988), .A1(N1678), .B0(N2420));
AOI21XL inst_cellmath__43_0_I1627 (.Y(N2596), .A0(N3045), .A1(N2670), .B0(N2621));
AOI21XL inst_cellmath__43_0_I1628 (.Y(N2346), .A0(N2802), .A1(N3388), .B0(N2372));
INVXL inst_cellmath__43_0_I1629 (.Y(N2093), .A(N2552));
INVXL inst_cellmath__43_0_I1630 (.Y(N2524), .A(N2120));
OAI21XL inst_cellmath__43_0_I1631 (.Y(N2950), .A0(N2093), .A1(N3095), .B0(N2524));
INVXL inst_cellmath__43_0_I1632 (.Y(N2698), .A(N2297));
INVXL inst_cellmath__43_0_I1633 (.Y(N3125), .A(N1868));
OAI21XL inst_cellmath__43_0_I1634 (.Y(N1595), .A0(N2698), .A1(N2025), .B0(N3125));
AOI21XL inst_cellmath__43_0_I1635 (.Y(N3305), .A0(N2045), .A1(N1562), .B0(N1621));
AOI21XL inst_cellmath__43_0_I1636 (.Y(N3053), .A0(N1795), .A1(N1777), .B0(N3332));
AOI21XL inst_cellmath__43_0_I1637 (.Y(N2809), .A0(N3509), .A1(N1992), .B0(N3077));
AOI21XL inst_cellmath__43_0_I1638 (.Y(N2558), .A0(N3260), .A1(N3490), .B0(N2832));
INVXL inst_cellmath__43_0_I1639 (.Y(N2303), .A(N3006));
INVXL inst_cellmath__43_0_I1640 (.Y(N2734), .A(N2584));
OAI21XL inst_cellmath__43_0_I1641 (.Y(N3160), .A0(N2303), .A1(N2423), .B0(N2734));
INVXL inst_cellmath__43_0_I1642 (.Y(N2908), .A(N2759));
INVXL inst_cellmath__43_0_I1643 (.Y(N3339), .A(N2330));
OAI21XL inst_cellmath__43_0_I1644 (.Y(N1802), .A0(N2908), .A1(N2135), .B0(N3339));
INVXL inst_cellmath__43_0_I1645 (.Y(N1552), .A(N2510));
INVXL inst_cellmath__43_0_I1646 (.Y(N1982), .A(N2078));
OAI21XL inst_cellmath__43_0_I1647 (.Y(N2410), .A0(N1552), .A1(N2848), .B0(N1982));
OR2XL inst_cellmath__43_0_I1648 (.Y(inst_cellmath__43[47]), .A(N2159), .B(N2741));
XNOR2X1 inst_cellmath__43_0_I1655 (.Y(inst_cellmath__43[23]), .A(N2845), .B(N2191));
XNOR2X1 inst_cellmath__43_0_I1656 (.Y(inst_cellmath__43[24]), .A(N2670), .B(N3045));
XOR2XL inst_cellmath__43_0_I1657 (.Y(inst_cellmath__43[25]), .A(N2596), .B(N1943));
XNOR2X1 inst_cellmath__43_0_I1658 (.Y(inst_cellmath__43[26]), .A(N3388), .B(N2802));
XOR2XL inst_cellmath__43_0_I1659 (.Y(inst_cellmath__43[27]), .A(N2346), .B(N1697));
XOR2XL inst_cellmath__43_0_I1660 (.Y(inst_cellmath__43[28]), .A(N3095), .B(N2552));
XNOR2X1 inst_cellmath__43_0_I1661 (.Y(inst_cellmath__43[29]), .A(N2950), .B(N3409));
XOR2XL inst_cellmath__43_0_I1662 (.Y(inst_cellmath__43[30]), .A(N2025), .B(N2297));
XNOR2X1 inst_cellmath__43_0_I1663 (.Y(inst_cellmath__43[31]), .A(N1595), .B(N3154));
XNOR2X1 inst_cellmath__43_0_I1664 (.Y(inst_cellmath__43[32]), .A(N1562), .B(N2045));
XOR2XL inst_cellmath__43_0_I1665 (.Y(inst_cellmath__43[33]), .A(N3305), .B(N2902));
XNOR2X1 inst_cellmath__43_0_I1666 (.Y(inst_cellmath__43[34]), .A(N1777), .B(N1795));
XOR2XL inst_cellmath__43_0_I1667 (.Y(inst_cellmath__43[35]), .A(N3053), .B(N2656));
XNOR2X1 inst_cellmath__43_0_I1668 (.Y(inst_cellmath__43[36]), .A(N1992), .B(N3509));
XOR2XL inst_cellmath__43_0_I1669 (.Y(inst_cellmath__43[37]), .A(N2809), .B(N2403));
XNOR2X1 inst_cellmath__43_0_I1670 (.Y(inst_cellmath__43[38]), .A(N3490), .B(N3260));
XOR2XL inst_cellmath__43_0_I1671 (.Y(inst_cellmath__43[39]), .A(N2558), .B(N2152));
XOR2XL inst_cellmath__43_0_I1672 (.Y(inst_cellmath__43[40]), .A(N2423), .B(N3006));
XNOR2X1 inst_cellmath__43_0_I1673 (.Y(inst_cellmath__43[41]), .A(N3160), .B(N1901));
XOR2XL inst_cellmath__43_0_I1674 (.Y(inst_cellmath__43[42]), .A(N2135), .B(N2759));
XNOR2X1 inst_cellmath__43_0_I1675 (.Y(inst_cellmath__43[43]), .A(N1802), .B(N1653));
XOR2XL inst_cellmath__43_0_I1676 (.Y(inst_cellmath__43[44]), .A(N2848), .B(N2510));
XNOR2X1 inst_cellmath__43_0_I1677 (.Y(inst_cellmath__43[45]), .A(N2410), .B(N3365));
XNOR2X1 inst_cellmath__43_0_I1678 (.Y(inst_cellmath__43[46]), .A(N2741), .B(N2159));
NOR2XL cynw_cm_float_mul_I1679 (.Y(N5430), .A(inst_cellmath__26), .B(inst_cellmath__22));
NOR2XL inst_cellmath__30__14__I1681 (.Y(N5437), .A(inst_cellmath__25), .B(inst_cellmath__21));
NAND2XL inst_cellmath__30__14__I1682 (.Y(N272), .A(N5437), .B(inst_cellmath__24));
OAI2BB1X1 cynw_cm_float_mul_I3432 (.Y(inst_cellmath__30), .A0N(N5430), .A1N(inst_cellmath__23), .B0(N272));
INVXL inst_cellmath__34_0_I1684 (.Y(N5452), .A(a_exp[7]));
XNOR2X1 inst_cellmath__34_0_I1685 (.Y(inst_cellmath__34[0]), .A(b_exp[0]), .B(a_exp[0]));
OR2XL inst_cellmath__34_0_I1686 (.Y(N5456), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 inst_cellmath__34_0_I1687 (.CO(N5449), .S(inst_cellmath__34[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(N5456));
ADDFX1 inst_cellmath__34_0_I1688 (.CO(N5468), .S(inst_cellmath__34[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(N5449));
ADDFX1 inst_cellmath__34_0_I1689 (.CO(N5480), .S(inst_cellmath__34[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(N5468));
ADDFX1 inst_cellmath__34_0_I1690 (.CO(N5462), .S(inst_cellmath__34[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(N5480));
ADDFX1 inst_cellmath__34_0_I1691 (.CO(N5477), .S(inst_cellmath__34[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(N5462));
ADDFX1 inst_cellmath__34_0_I1692 (.CO(N5457), .S(inst_cellmath__34[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(N5477));
ADDFX1 inst_cellmath__34_0_I1693 (.CO(N5472), .S(inst_cellmath__34[7]), .A(N5452), .B(b_exp[7]), .CI(N5457));
XNOR2X1 inst_cellmath__34_0_I1694 (.Y(inst_cellmath__34[8]), .A(a_exp[7]), .B(N5472));
NOR2XL inst_cellmath__34_0_I1695 (.Y(inst_cellmath__34[9]), .A(a_exp[7]), .B(N5472));
AND4XL inst_cellmath__41__24__I1696 (.Y(N5505), .A(inst_cellmath__34[0]), .B(inst_cellmath__34[1]), .C(inst_cellmath__34[2]), .D(inst_cellmath__34[3]));
NAND3XL inst_cellmath__41__24__I1697 (.Y(N5507), .A(inst_cellmath__34[4]), .B(inst_cellmath__34[7]), .C(inst_cellmath__34[5]));
NAND2XL inst_cellmath__41__24__I1698 (.Y(N5501), .A(inst_cellmath__34[6]), .B(N5505));
NOR2XL inst_cellmath__41__24__I1699 (.Y(N276), .A(N5507), .B(N5501));
NOR2XL andori2bb1_A_I3444 (.Y(N8078), .A(inst_cellmath__34[8]), .B(N276));
NOR2XL andori2bb1_A_I3445 (.Y(inst_cellmath__41), .A(N8078), .B(inst_cellmath__34[9]));
OR2XL cynw_cm_float_mul_I1702 (.Y(inst_cellmath__37), .A(inst_cellmath__30), .B(inst_cellmath__41));
NOR2XL inst_cellmath__35__16__I1703 (.Y(N5530), .A(inst_cellmath__34[0]), .B(inst_cellmath__34[9]));
NOR4BX1 inst_cellmath__35__16__I1704 (.Y(N5534), .AN(N5530), .B(inst_cellmath__34[1]), .C(inst_cellmath__34[8]), .D(inst_cellmath__34[2]));
NOR2XL inst_cellmath__35__16__I1705 (.Y(N5538), .A(inst_cellmath__34[7]), .B(inst_cellmath__34[6]));
OR3XL inst_cellmath__35__16__I1706 (.Y(N5529), .A(inst_cellmath__34[3]), .B(inst_cellmath__34[4]), .C(inst_cellmath__34[5]));
NAND3BXL inst_cellmath__35__16__I1707 (.Y(N273), .AN(N5529), .B(N5538), .C(N5534));
NOR3BXL cynw_cm_float_mul_I1708 (.Y(N269), .AN(inst_cellmath__25), .B(inst_cellmath__22), .C(inst_cellmath__24));
NOR3BXL cynw_cm_float_mul_I1709 (.Y(N270), .AN(inst_cellmath__26), .B(inst_cellmath__21), .C(inst_cellmath__23));
OR2XL cynw_cm_float_mul_I1710 (.Y(inst_cellmath__32), .A(N269), .B(N270));
NOR3XL inst_cellmath__60_0_I1711 (.Y(N5564), .A(inst_cellmath__32), .B(inst_cellmath__29), .C(inst_cellmath__34[9]));
NAND2XL inst_cellmath__60_0_I1712 (.Y(N5566), .A(N5564), .B(N273));
NOR2XL inst_cellmath__60_0_I1713 (.Y(inst_cellmath__60), .A(N5566), .B(inst_cellmath__37));
NAND3XL inst_cellmath__42__22__I3434 (.Y(N5580), .A(inst_cellmath__34[1]), .B(inst_cellmath__34[2]), .C(inst_cellmath__34[5]));
NAND4XL inst_cellmath__42__22__I3439 (.Y(N5575), .A(inst_cellmath__34[3]), .B(inst_cellmath__34[4]), .C(inst_cellmath__34[6]), .D(inst_cellmath__34[7]));
NOR2XL inst_cellmath__42__22__I1720 (.Y(N274), .A(N5580), .B(N5575));
NOR2XL andori2bb1_A_I3446 (.Y(N8085), .A(inst_cellmath__34[8]), .B(N274));
NOR2XL andori2bb1_A_I3447 (.Y(inst_cellmath__42), .A(N8085), .B(inst_cellmath__34[9]));
OR2XL cynw_cm_float_mul_I1723 (.Y(inst_cellmath__38), .A(inst_cellmath__30), .B(inst_cellmath__42));
NOR4X1 cynw_cm_float_mul_I1724 (.Y(inst_cellmath__61), .A(inst_cellmath__32), .B(inst_cellmath__29), .C(inst_cellmath__34[9]), .D(inst_cellmath__38));
MXI2XL cynw_cm_float_mul_I1725 (.Y(inst_cellmath__56), .A(inst_cellmath__60), .B(inst_cellmath__61), .S0(inst_cellmath__43[47]));
INVXL inst_cellmath__50_0_I1726 (.Y(inst_cellmath__50[0]), .A(inst_cellmath__34[0]));
NOR2BX1 inst_cellmath__50_0_I1727 (.Y(N5641), .AN(inst_cellmath__34[1]), .B(inst_cellmath__50[0]));
XNOR2X1 inst_cellmath__50_0_I1728 (.Y(inst_cellmath__50[1]), .A(inst_cellmath__50[0]), .B(inst_cellmath__34[1]));
NAND2XL inst_cellmath__50_0_I1729 (.Y(N5631), .A(inst_cellmath__34[2]), .B(N5641));
INVXL inst_cellmath__50_0_I1730 (.Y(N5622), .A(inst_cellmath__34[4]));
INVXL inst_cellmath__50_0_I1731 (.Y(N5633), .A(inst_cellmath__34[3]));
NOR3XL inst_cellmath__50_0_I1732 (.Y(N5620), .A(N5622), .B(N5633), .C(N5631));
NAND3XL inst_cellmath__50_0_I1733 (.Y(N5625), .A(inst_cellmath__34[5]), .B(N5620), .C(inst_cellmath__34[6]));
NAND2XL inst_cellmath__50_0_I1734 (.Y(N5627), .A(inst_cellmath__34[5]), .B(N5620));
XOR2XL inst_cellmath__50_0_I1735 (.Y(inst_cellmath__50[2]), .A(N5641), .B(inst_cellmath__34[2]));
XOR2XL inst_cellmath__50_0_I1736 (.Y(inst_cellmath__50[3]), .A(N5631), .B(N5633));
NOR2XL inst_cellmath__50_0_I1737 (.Y(N5618), .A(N5633), .B(N5631));
XNOR2X1 inst_cellmath__50_0_I1738 (.Y(inst_cellmath__50[4]), .A(N5622), .B(N5618));
XOR2XL inst_cellmath__50_0_I1739 (.Y(inst_cellmath__50[5]), .A(N5620), .B(inst_cellmath__34[5]));
XNOR2X1 inst_cellmath__50_0_I1740 (.Y(inst_cellmath__50[6]), .A(N5627), .B(inst_cellmath__34[6]));
XNOR2X1 inst_cellmath__50_0_I1741 (.Y(inst_cellmath__50[7]), .A(N5625), .B(inst_cellmath__34[7]));
OR3XL cynw_cm_float_mul_I1742 (.Y(inst_cellmath__54[7]), .A(inst_cellmath__29), .B(inst_cellmath__37), .C(inst_cellmath__38));
NOR2X1 inst_cellmath__64_2WWMM_I1744 (.Y(N5767), .A(inst_cellmath__43[47]), .B(inst_cellmath__56));
NOR2BX1 inst_cellmath__64_2WWMM_I1745 (.Y(N5682), .AN(inst_cellmath__43[47]), .B(inst_cellmath__56));
AOI22XL inst_cellmath__64_2WWMM_I1746 (.Y(N5694), .A0(inst_cellmath__50[0]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[0]));
AOI22XL inst_cellmath__64_2WWMM_I1747 (.Y(N5743), .A0(inst_cellmath__50[1]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[1]));
AOI22XL inst_cellmath__64_2WWMM_I1748 (.Y(N5680), .A0(inst_cellmath__50[2]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[2]));
AOI22XL inst_cellmath__64_2WWMM_I1749 (.Y(N5729), .A0(inst_cellmath__50[3]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[3]));
AOI22XL inst_cellmath__64_2WWMM_I1750 (.Y(N5778), .A0(inst_cellmath__50[4]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[4]));
AOI22XL inst_cellmath__64_2WWMM_I1751 (.Y(N5714), .A0(inst_cellmath__50[5]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[5]));
AOI22XL inst_cellmath__64_2WWMM_I1752 (.Y(N5762), .A0(inst_cellmath__50[6]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[6]));
AOI22XL inst_cellmath__64_2WWMM_I1753 (.Y(N5700), .A0(inst_cellmath__50[7]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__34[7]));
AOI22XL inst_cellmath__64_2WWMM_I1754 (.Y(N5750), .A0(inst_cellmath__43[24]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[23]));
AOI22XL inst_cellmath__64_2WWMM_I1755 (.Y(N5687), .A0(inst_cellmath__43[25]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[24]));
AOI22XL inst_cellmath__64_2WWMM_I1756 (.Y(N5735), .A0(inst_cellmath__43[26]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[25]));
AOI22XL inst_cellmath__64_2WWMM_I1757 (.Y(N5672), .A0(inst_cellmath__43[27]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[26]));
AOI22XL inst_cellmath__64_2WWMM_I1758 (.Y(N5722), .A0(inst_cellmath__43[28]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[27]));
AOI22XL inst_cellmath__64_2WWMM_I1759 (.Y(N5770), .A0(inst_cellmath__43[29]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[28]));
AOI22XL inst_cellmath__64_2WWMM_I1760 (.Y(N5707), .A0(inst_cellmath__43[30]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[29]));
AOI22XL inst_cellmath__64_2WWMM_I1761 (.Y(N5755), .A0(inst_cellmath__43[31]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[30]));
AOI22XL inst_cellmath__64_2WWMM_I1762 (.Y(N5692), .A0(inst_cellmath__43[32]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[31]));
AOI22XL inst_cellmath__64_2WWMM_I1763 (.Y(N5741), .A0(inst_cellmath__43[33]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[32]));
AOI22XL inst_cellmath__64_2WWMM_I1764 (.Y(N5677), .A0(inst_cellmath__43[34]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[33]));
AOI22XL inst_cellmath__64_2WWMM_I1765 (.Y(N5727), .A0(inst_cellmath__43[35]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[34]));
AOI22XL inst_cellmath__64_2WWMM_I1766 (.Y(N5776), .A0(inst_cellmath__43[36]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[35]));
AOI22XL inst_cellmath__64_2WWMM_I1767 (.Y(N5711), .A0(inst_cellmath__43[37]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[36]));
AOI22XL inst_cellmath__64_2WWMM_I1768 (.Y(N5759), .A0(inst_cellmath__43[38]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[37]));
AOI22XL inst_cellmath__64_2WWMM_I1769 (.Y(N5697), .A0(inst_cellmath__43[39]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[38]));
AOI22XL inst_cellmath__64_2WWMM_I1770 (.Y(N5747), .A0(inst_cellmath__43[40]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[39]));
AOI22XL inst_cellmath__64_2WWMM_I1771 (.Y(N5684), .A0(inst_cellmath__43[41]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[40]));
AOI22XL inst_cellmath__64_2WWMM_I1772 (.Y(N5732), .A0(inst_cellmath__43[42]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[41]));
AOI22XL inst_cellmath__64_2WWMM_I1773 (.Y(N5669), .A0(inst_cellmath__43[43]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[42]));
AOI22XL inst_cellmath__64_2WWMM_I1774 (.Y(N5719), .A0(inst_cellmath__43[44]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[43]));
AOI22XL inst_cellmath__64_2WWMM_I1775 (.Y(N5766), .A0(inst_cellmath__43[45]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[44]));
AOI22XL inst_cellmath__64_2WWMM_I1776 (.Y(N5705), .A0(inst_cellmath__43[46]), .A1(N5682), .B0(N5767), .B1(inst_cellmath__43[45]));
NAND2XL inst_cellmath__64_2WWMM_I1777 (.Y(N5701), .A(inst_cellmath__56), .B(inst_cellmath__54[7]));
NAND2X1 inst_cellmath__64_2WWMM_I1778 (.Y(N5673), .A(inst_cellmath__56), .B(inst_cellmath__29));
NAND2XL inst_cellmath__64_2WWMM_I1779 (.Y(x[23]), .A(N5701), .B(N5694));
NAND2XL inst_cellmath__64_2WWMM_I1780 (.Y(x[24]), .A(N5701), .B(N5743));
NAND2XL inst_cellmath__64_2WWMM_I1781 (.Y(x[25]), .A(N5701), .B(N5680));
NAND2XL inst_cellmath__64_2WWMM_I1782 (.Y(x[26]), .A(N5701), .B(N5729));
NAND2XL inst_cellmath__64_2WWMM_I1783 (.Y(x[27]), .A(N5701), .B(N5778));
NAND2XL inst_cellmath__64_2WWMM_I1784 (.Y(x[28]), .A(N5701), .B(N5714));
NAND2XL inst_cellmath__64_2WWMM_I1785 (.Y(x[29]), .A(N5701), .B(N5762));
OAI2BB1X1 inst_cellmath__64_2WWMM_I1786 (.Y(x[30]), .A0N(inst_cellmath__56), .A1N(inst_cellmath__54[7]), .B0(N5700));
NAND2XL inst_cellmath__64_2WWMM_I1787 (.Y(x[0]), .A(N5673), .B(N5750));
NAND2XL inst_cellmath__64_2WWMM_I1788 (.Y(x[1]), .A(N5673), .B(N5687));
NAND2XL inst_cellmath__64_2WWMM_I1789 (.Y(x[2]), .A(N5673), .B(N5735));
NAND2XL inst_cellmath__64_2WWMM_I1790 (.Y(x[3]), .A(N5673), .B(N5672));
NAND2XL inst_cellmath__64_2WWMM_I1791 (.Y(x[4]), .A(N5673), .B(N5722));
NAND2XL inst_cellmath__64_2WWMM_I1792 (.Y(x[5]), .A(N5673), .B(N5770));
NAND2XL inst_cellmath__64_2WWMM_I1793 (.Y(x[6]), .A(N5673), .B(N5707));
NAND2XL inst_cellmath__64_2WWMM_I1794 (.Y(x[7]), .A(N5673), .B(N5755));
NAND2XL inst_cellmath__64_2WWMM_I1795 (.Y(x[8]), .A(N5673), .B(N5692));
NAND2XL inst_cellmath__64_2WWMM_I1796 (.Y(x[9]), .A(N5673), .B(N5741));
NAND2XL inst_cellmath__64_2WWMM_I1797 (.Y(x[10]), .A(N5673), .B(N5677));
NAND2XL inst_cellmath__64_2WWMM_I1798 (.Y(x[11]), .A(N5673), .B(N5727));
NAND2XL inst_cellmath__64_2WWMM_I1799 (.Y(x[12]), .A(N5673), .B(N5776));
NAND2XL inst_cellmath__64_2WWMM_I1800 (.Y(x[13]), .A(N5673), .B(N5711));
NAND2XL inst_cellmath__64_2WWMM_I1801 (.Y(x[14]), .A(N5673), .B(N5759));
NAND2XL inst_cellmath__64_2WWMM_I1802 (.Y(x[15]), .A(N5673), .B(N5697));
NAND2XL inst_cellmath__64_2WWMM_I1803 (.Y(x[16]), .A(N5673), .B(N5747));
NAND2XL inst_cellmath__64_2WWMM_I1804 (.Y(x[17]), .A(N5673), .B(N5684));
NAND2XL inst_cellmath__64_2WWMM_I1805 (.Y(x[18]), .A(N5673), .B(N5732));
NAND2XL inst_cellmath__64_2WWMM_I1806 (.Y(x[19]), .A(N5673), .B(N5669));
NAND2XL inst_cellmath__64_2WWMM_I1807 (.Y(x[20]), .A(N5673), .B(N5719));
NAND2XL inst_cellmath__64_2WWMM_I1808 (.Y(x[21]), .A(N5673), .B(N5766));
NAND2XL inst_cellmath__64_2WWMM_I1809 (.Y(x[22]), .A(N5673), .B(N5705));
assign inst_cellmath__43[0] = 1'B0;
assign inst_cellmath__43[1] = 1'B0;
assign inst_cellmath__43[2] = 1'B0;
assign inst_cellmath__43[3] = 1'B0;
assign inst_cellmath__43[4] = 1'B0;
assign inst_cellmath__43[5] = 1'B0;
assign inst_cellmath__43[6] = 1'B0;
assign inst_cellmath__43[7] = 1'B0;
assign inst_cellmath__43[8] = 1'B0;
assign inst_cellmath__43[9] = 1'B0;
assign inst_cellmath__43[10] = 1'B0;
assign inst_cellmath__43[11] = 1'B0;
assign inst_cellmath__43[12] = 1'B0;
assign inst_cellmath__43[13] = 1'B0;
assign inst_cellmath__43[14] = 1'B0;
assign inst_cellmath__43[15] = 1'B0;
assign inst_cellmath__43[16] = 1'B0;
assign inst_cellmath__43[17] = 1'B0;
assign inst_cellmath__43[18] = 1'B0;
assign inst_cellmath__43[19] = 1'B0;
assign inst_cellmath__43[20] = 1'B0;
assign inst_cellmath__43[21] = 1'B0;
assign inst_cellmath__43[22] = 1'B0;
assign inst_cellmath__54[0] = 1'B0;
assign inst_cellmath__54[1] = 1'B0;
assign inst_cellmath__54[2] = 1'B0;
assign inst_cellmath__54[3] = 1'B0;
assign inst_cellmath__54[4] = 1'B0;
assign inst_cellmath__54[5] = 1'B0;
assign inst_cellmath__54[6] = 1'B0;
endmodule

/* CADENCE  urX3SwHXrh8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



