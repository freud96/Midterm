/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:23:43 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24;
wire [8:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42;
wire [22:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82;
wire [0:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1;
wire [29:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195;
wire [32:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198;
wire [49:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201;
wire [46:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1;
wire [30:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210;
wire [4:0] DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215;
wire  DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712,
	DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720;
wire N9100,N18660,N18664,N18667,N18678,N18835,N18839 
	,N18879,N18881,N18886,N18971,N18990,N19000,N19010,N19020 
	,N19030,N19040,N19050,N19060,N19070,N19080,N19099,N19109 
	,N19119,N19129,N19139,N19149,N19159,N19223,N19233,N19275 
	,N19410,N19633,N19768,N19891,N19900,N19909,N20144,N20175 
	,N20182,N20492,N20538,N20660,N21070,N21075,N21080,N21085 
	,N21090,N21100,N21105,N21765,N21769,N21782,N21795,N21988 
	,N21993,N21999,N22003,N22305,N22309,N22618,N22929,N22939 
	,N22949,N22959,N22969,N22979,N22989,N23008,N23018,N23035 
	,N23050,N23060,N23070,N23080,N23090,N23100,N23110,N23120 
	,N23130,N23140,N23142,N23333,N23335,N23378,N23556,N23579 
	,N23859,N23861,N23943,N23945,N24239,N24241,N24248,N24250 
	,N24268,N24432,N24633,N24635,N24642,N24644,N24653,N24662 
	,N25288,N25295,N25297,N25313,N25457,N25627,N25766,N25768 
	,N25852,N25854,N26198,N26206,N26208,N26228,N26230,N26236 
	,N26238,N26244,N26246,N26248,N26252,N26254,N26256,N26646 
	,N26654,N26704,N26726,N26734,N26736,N26742,N26744,N26750 
	,N26752,N26758,N26760,N26766,N26768,N27092,N27094,N27100 
	,N27102,N27231,N27448,N27456,N27640,N27844,N27939,N28088 
	,N28113,N28287,N28313,N29392,N29396,N29398,N29426,N29430 
	,N29442,N29446,N29448,N29450,N29452,N29454,N29456,N29458 
	,N29460,N29462,N29464,N29466,N29468,N29470,N29472,N29474 
	,N29476,N29478,N29480,N29482,N29484,N29486,N29488,N29490 
	,N29492,N29494,N29496,N29498,N29502,N29506,N29510,N29556 
	,N29560,N29566,N29570,N29580,N29592,N29598,N29610,N29612 
	,N29614,N29616,N29618,N29620,N29622,N29624,N29626,N29653 
	,N29655,N29667,N29669,N29673,N29679,N29681,N30223,N30224 
	,N30225,N30226,N30227,N30228,N30229,N30230,N30231,N30232 
	,N30233,N30234,N30235,N30236,N30237,N30238,N30239,N30240 
	,N30241,N30242,N30243,N30244,N30245,N30246,N30247,N30248 
	,N30249,N30250,N30251,N30252,N30253,N30254,N30255,N30256 
	,N30257,N30258,N30259,N30260,N30261,N30262,N30263,N30264 
	,N30265,N30266,N30267,N30268,N30269,N30270,N30271,N30272 
	,N30273,N30274,N30275,N30276,N30277,N30278,N30279,N30280 
	,N30281,N30282,N30283,N30284,N30285,N30286,N30287,N30288 
	,N30289,N30290,N30291,N30292,N30293,N30294,N30295,N30296 
	,N30297,N30298,N30299,N30300,N30301,N30302,N30303,N30304 
	,N30305,N30306,N30307,N30308,N30309,N30310,N30311,N30312 
	,N30313,N30315,N30316,N30323,N30329,N30336,N30343,N30352 
	,N30360,N30368,N30373;
reg x_reg_L0_31__retimed_I15390_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15390_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002;
	end
assign N29681 = x_reg_L0_31__retimed_I15390_QOUT;
reg x_reg_L0_31__retimed_I15389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15389_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921;
	end
assign N29679 = x_reg_L0_31__retimed_I15389_QOUT;
reg x_reg_L0_31__retimed_I15387_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15387_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330;
	end
assign N29673 = x_reg_L0_31__retimed_I15387_QOUT;
reg x_reg_L0_31__retimed_I15386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15386_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355;
	end
assign N29669 = x_reg_L0_31__retimed_I15386_QOUT;
reg x_reg_L0_31__retimed_I15385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15385_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276;
	end
assign N29667 = x_reg_L0_31__retimed_I15385_QOUT;
reg x_reg_L0_31__retimed_I15380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15380_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109;
	end
assign N29655 = x_reg_L0_31__retimed_I15380_QOUT;
reg x_reg_L0_31__retimed_I15379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15379_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746;
	end
assign N29653 = x_reg_L0_31__retimed_I15379_QOUT;
reg x_reg_L0_31__retimed_I15368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15368_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486;
	end
assign N29626 = x_reg_L0_31__retimed_I15368_QOUT;
reg x_reg_L0_31__retimed_I15367_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15367_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098;
	end
assign N29624 = x_reg_L0_31__retimed_I15367_QOUT;
reg x_reg_L0_31__retimed_I15366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15366_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668;
	end
assign N29622 = x_reg_L0_31__retimed_I15366_QOUT;
reg x_reg_L0_31__retimed_I15365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15365_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982;
	end
assign N29620 = x_reg_L0_31__retimed_I15365_QOUT;
reg x_reg_L0_31__retimed_I15364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15364_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147;
	end
assign N29618 = x_reg_L0_31__retimed_I15364_QOUT;
reg x_reg_L0_31__retimed_I15363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15363_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791;
	end
assign N29616 = x_reg_L0_31__retimed_I15363_QOUT;
reg x_reg_L0_31__retimed_I15362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15362_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[32];
	end
assign N29614 = x_reg_L0_31__retimed_I15362_QOUT;
reg x_reg_L0_31__retimed_I15361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15361_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601;
	end
assign N29612 = x_reg_L0_31__retimed_I15361_QOUT;
reg x_reg_L0_31__retimed_I15360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15360_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212;
	end
assign N29610 = x_reg_L0_31__retimed_I15360_QOUT;
reg x_reg_L0_31__retimed_I15354_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15354_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[31];
	end
assign N29598 = x_reg_L0_31__retimed_I15354_QOUT;
reg x_reg_L0_31__retimed_I15351_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15351_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[30];
	end
assign N29592 = x_reg_L0_31__retimed_I15351_QOUT;
reg x_reg_L0_31__retimed_I15345_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15345_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[29];
	end
assign N29580 = x_reg_L0_31__retimed_I15345_QOUT;
reg x_reg_L0_31__retimed_I15340_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15340_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[27];
	end
assign N29570 = x_reg_L0_31__retimed_I15340_QOUT;
reg x_reg_L0_31__retimed_I15338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15338_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918;
	end
assign N29566 = x_reg_L0_31__retimed_I15338_QOUT;
reg x_reg_L0_31__retimed_I15335_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15335_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[26];
	end
assign N29560 = x_reg_L0_31__retimed_I15335_QOUT;
reg x_reg_L0_31__retimed_I15333_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15333_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153;
	end
assign N29556 = x_reg_L0_31__retimed_I15333_QOUT;
assign N30223 = !N29556;
assign N30224 = !N30223;
reg x_reg_L0_31__retimed_I15310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15310_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415;
	end
assign N29510 = x_reg_L0_31__retimed_I15310_QOUT;
reg x_reg_L0_31__retimed_I15308_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15308_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222;
	end
assign N29506 = x_reg_L0_31__retimed_I15308_QOUT;
reg x_reg_L0_31__retimed_I15306_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15306_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080;
	end
assign N29502 = x_reg_L0_31__retimed_I15306_QOUT;
reg x_reg_L0_31__retimed_I15304_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15304_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890;
	end
assign N29498 = x_reg_L0_31__retimed_I15304_QOUT;
reg x_reg_L0_31__retimed_I15303_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15303_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089;
	end
assign N29496 = x_reg_L0_31__retimed_I15303_QOUT;
reg x_reg_L0_31__retimed_I15302_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15302_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744;
	end
assign N29494 = x_reg_L0_31__retimed_I15302_QOUT;
reg x_reg_L0_31__retimed_I15301_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15301_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983;
	end
assign N29492 = x_reg_L0_31__retimed_I15301_QOUT;
reg x_reg_L0_31__retimed_I15300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15300_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611;
	end
assign N29490 = x_reg_L0_31__retimed_I15300_QOUT;
reg x_reg_L0_31__retimed_I15299_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15299_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072;
	end
assign N29488 = x_reg_L0_31__retimed_I15299_QOUT;
reg x_reg_L0_31__retimed_I15298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15298_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731;
	end
assign N29486 = x_reg_L0_31__retimed_I15298_QOUT;
reg x_reg_L0_31__retimed_I15297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15297_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860;
	end
assign N29484 = x_reg_L0_31__retimed_I15297_QOUT;
reg x_reg_L0_31__retimed_I15296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15296_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469;
	end
assign N29482 = x_reg_L0_31__retimed_I15296_QOUT;
reg x_reg_L0_31__retimed_I15295_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15295_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237;
	end
assign N29480 = x_reg_L0_31__retimed_I15295_QOUT;
reg x_reg_L0_31__retimed_I15294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15294_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866;
	end
assign N29478 = x_reg_L0_31__retimed_I15294_QOUT;
reg x_reg_L0_31__retimed_I15293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15293_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120;
	end
assign N29476 = x_reg_L0_31__retimed_I15293_QOUT;
reg x_reg_L0_31__retimed_I15292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15292_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771;
	end
assign N29474 = x_reg_L0_31__retimed_I15292_QOUT;
reg x_reg_L0_31__retimed_I15291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15291_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417;
	end
assign N29472 = x_reg_L0_31__retimed_I15291_QOUT;
reg x_reg_L0_31__retimed_I15290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15290_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035;
	end
assign N29470 = x_reg_L0_31__retimed_I15290_QOUT;
reg x_reg_L0_31__retimed_I15289_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15289_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167;
	end
assign N29468 = x_reg_L0_31__retimed_I15289_QOUT;
reg x_reg_L0_31__retimed_I15288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15288_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807;
	end
assign N29466 = x_reg_L0_31__retimed_I15288_QOUT;
reg x_reg_L0_31__retimed_I15287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15287_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202;
	end
assign N29464 = x_reg_L0_31__retimed_I15287_QOUT;
reg x_reg_L0_31__retimed_I15286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15286_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846;
	end
assign N29462 = x_reg_L0_31__retimed_I15286_QOUT;
reg x_reg_L0_31__retimed_I15285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15285_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497;
	end
assign N29460 = x_reg_L0_31__retimed_I15285_QOUT;
reg x_reg_L0_31__retimed_I15284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15284_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105;
	end
assign N29458 = x_reg_L0_31__retimed_I15284_QOUT;
reg x_reg_L0_31__retimed_I15283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15283_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156;
	end
assign N29456 = x_reg_L0_31__retimed_I15283_QOUT;
reg x_reg_L0_31__retimed_I15282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15282_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798;
	end
assign N29454 = x_reg_L0_31__retimed_I15282_QOUT;
reg x_reg_L0_31__retimed_I15281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15281_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789;
	end
assign N29452 = x_reg_L0_31__retimed_I15281_QOUT;
reg x_reg_L0_31__retimed_I15280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15280_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124;
	end
assign N29450 = x_reg_L0_31__retimed_I15280_QOUT;
reg x_reg_L0_31__retimed_I15279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15279_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811;
	end
assign N29448 = x_reg_L0_31__retimed_I15279_QOUT;
reg x_reg_L0_31__retimed_I15278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15278_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426;
	end
assign N29446 = x_reg_L0_31__retimed_I15278_QOUT;
reg x_reg_L0_31__retimed_I15276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15276_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[24];
	end
assign N29442 = x_reg_L0_31__retimed_I15276_QOUT;
reg x_reg_L0_31__retimed_I15270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15270_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[25];
	end
assign N29430 = x_reg_L0_31__retimed_I15270_QOUT;
reg x_reg_L0_31__retimed_I15268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15268_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[28];
	end
assign N29426 = x_reg_L0_31__retimed_I15268_QOUT;
reg x_reg_L0_31__retimed_I15255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15255_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397;
	end
assign N29398 = x_reg_L0_31__retimed_I15255_QOUT;
reg x_reg_L0_31__retimed_I15254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15254_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015;
	end
assign N29396 = x_reg_L0_31__retimed_I15254_QOUT;
reg x_reg_L0_31__retimed_I15252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I15252_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[22];
	end
assign N29392 = x_reg_L0_31__retimed_I15252_QOUT;
reg x_reg_L0_31__retimed_I14964_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14964_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[18];
	end
assign N28313 = x_reg_L0_31__retimed_I14964_QOUT;
reg x_reg_L0_31__retimed_I14962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14962_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20];
	end
assign N28287 = x_reg_L0_31__retimed_I14962_QOUT;
reg x_reg_L0_31__retimed_I14921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14921_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19];
	end
assign N28113 = x_reg_L0_31__retimed_I14921_QOUT;
assign N30225 = !N28113;
assign N30226 = !N30225;
reg x_reg_L0_31__retimed_I14912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14912_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21];
	end
assign N28088 = x_reg_L0_31__retimed_I14912_QOUT;
reg x_reg_L0_31__retimed_I14868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14868_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[23];
	end
assign N27939 = x_reg_L0_31__retimed_I14868_QOUT;
reg x_reg_L0_31__retimed_I14846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14846_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564;
	end
assign N27844 = x_reg_L0_31__retimed_I14846_QOUT;
reg x_reg_L0_31__retimed_I14791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14791_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476;
	end
assign N27640 = x_reg_L0_31__retimed_I14791_QOUT;
reg x_reg_L0_31__retimed_I14734_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14734_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344;
	end
assign N27456 = x_reg_L0_31__retimed_I14734_QOUT;
reg x_reg_L0_31__retimed_I14731_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14731_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030;
	end
assign N27448 = x_reg_L0_31__retimed_I14731_QOUT;
reg x_reg_L0_31__retimed_I14653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14653_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717;
	end
assign N27231 = x_reg_L0_31__retimed_I14653_QOUT;
reg x_reg_L0_31__retimed_I14604_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14604_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857;
	end
assign N27102 = x_reg_L0_31__retimed_I14604_QOUT;
reg x_reg_L0_31__retimed_I14603_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14603_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840;
	end
assign N27100 = x_reg_L0_31__retimed_I14603_QOUT;
reg x_reg_L0_31__retimed_I14601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14601_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872;
	end
assign N27094 = x_reg_L0_31__retimed_I14601_QOUT;
reg x_reg_L0_31__retimed_I14600_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14600_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127;
	end
assign N27092 = x_reg_L0_31__retimed_I14600_QOUT;
reg x_reg_L0_31__retimed_I14504_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14504_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039;
	end
assign N26768 = x_reg_L0_31__retimed_I14504_QOUT;
reg x_reg_L0_31__retimed_I14503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14503_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021;
	end
assign N26766 = x_reg_L0_31__retimed_I14503_QOUT;
reg x_reg_L0_31__retimed_I14501_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14501_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739;
	end
assign N26760 = x_reg_L0_31__retimed_I14501_QOUT;
reg x_reg_L0_31__retimed_I14500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14500_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134;
	end
assign N26758 = x_reg_L0_31__retimed_I14500_QOUT;
reg x_reg_L0_31__retimed_I14498_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14498_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073;
	end
assign N26752 = x_reg_L0_31__retimed_I14498_QOUT;
reg x_reg_L0_31__retimed_I14497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14497_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758;
	end
assign N26750 = x_reg_L0_31__retimed_I14497_QOUT;
reg x_reg_L0_31__retimed_I14495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14495_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364;
	end
assign N26744 = x_reg_L0_31__retimed_I14495_QOUT;
reg x_reg_L0_31__retimed_I14494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14494_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108;
	end
assign N26742 = x_reg_L0_31__retimed_I14494_QOUT;
reg x_reg_L0_31__retimed_I14492_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14492_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760;
	end
assign N26736 = x_reg_L0_31__retimed_I14492_QOUT;
reg x_reg_L0_31__retimed_I14491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14491_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243;
	end
assign N26734 = x_reg_L0_31__retimed_I14491_QOUT;
reg x_reg_L0_31__retimed_I14488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14488_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757;
	end
assign N26726 = x_reg_L0_31__retimed_I14488_QOUT;
reg x_reg_L0_31__retimed_I14479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14479_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092;
	end
assign N26704 = x_reg_L0_31__retimed_I14479_QOUT;
reg x_reg_L0_31__retimed_I14458_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14458_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773;
	end
assign N26654 = x_reg_L0_31__retimed_I14458_QOUT;
reg x_reg_L0_31__retimed_I14455_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14455_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227;
	end
assign N26646 = x_reg_L0_31__retimed_I14455_QOUT;
reg x_reg_L0_31__retimed_I14320_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14320_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156;
	end
assign N26256 = x_reg_L0_31__retimed_I14320_QOUT;
reg x_reg_L0_31__retimed_I14319_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14319_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408;
	end
assign N26254 = x_reg_L0_31__retimed_I14319_QOUT;
reg x_reg_L0_31__retimed_I14318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14318_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607;
	end
assign N26252 = x_reg_L0_31__retimed_I14318_QOUT;
reg x_reg_L0_31__retimed_I14317_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14317_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026;
	end
assign N26248 = x_reg_L0_31__retimed_I14317_QOUT;
reg x_reg_L0_31__retimed_I14316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14316_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265;
	end
assign N26246 = x_reg_L0_31__retimed_I14316_QOUT;
reg x_reg_L0_31__retimed_I14315_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14315_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208;
	end
assign N26244 = x_reg_L0_31__retimed_I14315_QOUT;
reg x_reg_L0_31__retimed_I14313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14313_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903;
	end
assign N26238 = x_reg_L0_31__retimed_I14313_QOUT;
reg x_reg_L0_31__retimed_I14312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14312_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085;
	end
assign N26236 = x_reg_L0_31__retimed_I14312_QOUT;
reg x_reg_L0_31__retimed_I14310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14310_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816;
	end
assign N26230 = x_reg_L0_31__retimed_I14310_QOUT;
reg x_reg_L0_31__retimed_I14309_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14309_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370;
	end
assign N26228 = x_reg_L0_31__retimed_I14309_QOUT;
reg x_reg_L0_31__retimed_I14301_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14301_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035;
	end
assign N26208 = x_reg_L0_31__retimed_I14301_QOUT;
reg x_reg_L0_31__retimed_I14300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14300_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852;
	end
assign N26206 = x_reg_L0_31__retimed_I14300_QOUT;
reg x_reg_L0_31__retimed_I14297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14297_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742;
	end
assign N26198 = x_reg_L0_31__retimed_I14297_QOUT;
reg x_reg_L0_31__retimed_I14154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14154_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310;
	end
assign N25854 = x_reg_L0_31__retimed_I14154_QOUT;
assign N30227 = !N25854;
assign N30228 = !N30227;
reg x_reg_L0_31__retimed_I14153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14153_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975;
	end
assign N25852 = x_reg_L0_31__retimed_I14153_QOUT;
assign N30229 = !N25852;
assign N30230 = !N30229;
reg x_reg_L0_31__retimed_I14121_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14121_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710;
	end
assign N25768 = x_reg_L0_31__retimed_I14121_QOUT;
reg x_reg_L0_31__retimed_I14120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14120_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687;
	end
assign N25766 = x_reg_L0_31__retimed_I14120_QOUT;
reg x_reg_L0_31__retimed_I14062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I14062_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666;
	end
assign N25627 = x_reg_L0_31__retimed_I14062_QOUT;
reg x_reg_L0_31__retimed_I13990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13990_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219;
	end
assign N25457 = x_reg_L0_31__retimed_I13990_QOUT;
assign N30231 = !N25457;
assign N30232 = !N30231;
reg x_reg_L0_31__retimed_I13930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13930_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108;
	end
assign N25313 = x_reg_L0_31__retimed_I13930_QOUT;
assign N30233 = !N25313;
assign N30234 = !N30233;
reg x_reg_L0_31__retimed_I13923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13923_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352;
	end
assign N25297 = x_reg_L0_31__retimed_I13923_QOUT;
assign N30235 = !N25297;
assign N30236 = !N30235;
reg x_reg_L0_31__retimed_I13922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13922_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745;
	end
assign N25295 = x_reg_L0_31__retimed_I13922_QOUT;
assign N30237 = !N25295;
assign N30238 = !N30237;
reg x_reg_L0_31__retimed_I13919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13919_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774;
	end
assign N25288 = x_reg_L0_31__retimed_I13919_QOUT;
assign N30239 = !N25288;
assign N30240 = !N30239;
reg x_reg_L0_31__retimed_I13661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13661_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894;
	end
assign N24662 = x_reg_L0_31__retimed_I13661_QOUT;
assign N30241 = !N24662;
assign N30242 = !N30241;
reg x_reg_L0_31__retimed_I13657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13657_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284;
	end
assign N24653 = x_reg_L0_31__retimed_I13657_QOUT;
assign N30243 = !N24653;
assign N30244 = !N30243;
reg x_reg_L0_31__retimed_I13653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13653_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125;
	end
assign N24644 = x_reg_L0_31__retimed_I13653_QOUT;
assign N30245 = !N24644;
assign N30246 = !N30245;
reg x_reg_L0_31__retimed_I13652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13652_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517;
	end
assign N24642 = x_reg_L0_31__retimed_I13652_QOUT;
assign N30247 = !N24642;
assign N30248 = !N30247;
reg x_reg_L0_31__retimed_I13649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13649_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255;
	end
assign N24635 = x_reg_L0_31__retimed_I13649_QOUT;
assign N30249 = !N24635;
assign N30250 = !N30249;
reg x_reg_L0_31__retimed_I13648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13648_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914;
	end
assign N24633 = x_reg_L0_31__retimed_I13648_QOUT;
assign N30251 = !N24633;
assign N30252 = !N30251;
reg x_reg_L0_31__retimed_I13572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13572_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852;
	end
assign N24432 = x_reg_L0_31__retimed_I13572_QOUT;
reg x_reg_L0_31__retimed_I13503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13503_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677;
	end
assign N24268 = x_reg_L0_31__retimed_I13503_QOUT;
assign N30253 = !N24268;
assign N30254 = !N30253;
reg x_reg_L0_31__retimed_I13495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13495_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044;
	end
assign N24250 = x_reg_L0_31__retimed_I13495_QOUT;
assign N30255 = !N24250;
assign N30256 = !N30255;
reg x_reg_L0_31__retimed_I13494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13494_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236;
	end
assign N24248 = x_reg_L0_31__retimed_I13494_QOUT;
assign N30257 = !N24248;
assign N30258 = !N30257;
reg x_reg_L0_31__retimed_I13491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13491_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064;
	end
assign N24241 = x_reg_L0_31__retimed_I13491_QOUT;
assign N30259 = !N24241;
assign N30260 = !N30259;
reg x_reg_L0_31__retimed_I13490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13490_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447;
	end
assign N24239 = x_reg_L0_31__retimed_I13490_QOUT;
assign N30261 = !N24239;
assign N30262 = !N30261;
reg x_reg_L0_31__retimed_I13379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13379_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821;
	end
assign N23945 = x_reg_L0_31__retimed_I13379_QOUT;
reg x_reg_L0_31__retimed_I13378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13378_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073;
	end
assign N23943 = x_reg_L0_31__retimed_I13378_QOUT;
reg x_reg_L0_31__retimed_I13344_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13344_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832;
	end
assign N23861 = x_reg_L0_31__retimed_I13344_QOUT;
assign N30263 = !N23861;
assign N30264 = !N30263;
reg x_reg_L0_31__retimed_I13343_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13343_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191;
	end
assign N23859 = x_reg_L0_31__retimed_I13343_QOUT;
assign N30265 = !N23859;
assign N30266 = !N30265;
reg x_reg_L0_31__retimed_I13240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13240_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181;
	end
assign N23579 = x_reg_L0_31__retimed_I13240_QOUT;
reg x_reg_L0_31__retimed_I13231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13231_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851;
	end
assign N23556 = x_reg_L0_31__retimed_I13231_QOUT;
assign N30267 = !N23556;
assign N30268 = !N30267;
reg x_reg_L0_31__retimed_I13163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13163_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[0];
	end
assign N23378 = x_reg_L0_31__retimed_I13163_QOUT;
reg x_reg_L0_31__retimed_I13148_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13148_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763;
	end
assign N23335 = x_reg_L0_31__retimed_I13148_QOUT;
reg x_reg_L0_31__retimed_I13147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13147_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844;
	end
assign N23333 = x_reg_L0_31__retimed_I13147_QOUT;
reg x_reg_L0_31__retimed_I13074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13074_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[38];
	end
assign N23142 = x_reg_L0_31__retimed_I13074_QOUT;
reg x_reg_L0_31__retimed_I13073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13073_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[20];
	end
assign N23140 = x_reg_L0_31__retimed_I13073_QOUT;
reg x_reg_L0_31__retimed_I13070_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13070_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[19];
	end
assign N23130 = x_reg_L0_31__retimed_I13070_QOUT;
reg x_reg_L0_31__retimed_I13067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13067_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[18];
	end
assign N23120 = x_reg_L0_31__retimed_I13067_QOUT;
reg x_reg_L0_31__retimed_I13064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13064_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[17];
	end
assign N23110 = x_reg_L0_31__retimed_I13064_QOUT;
reg x_reg_L0_31__retimed_I13061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13061_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[16];
	end
assign N23100 = x_reg_L0_31__retimed_I13061_QOUT;
reg x_reg_L0_31__retimed_I13058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13058_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[15];
	end
assign N23090 = x_reg_L0_31__retimed_I13058_QOUT;
reg x_reg_L0_31__retimed_I13055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13055_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[14];
	end
assign N23080 = x_reg_L0_31__retimed_I13055_QOUT;
reg x_reg_L0_31__retimed_I13052_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13052_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[13];
	end
assign N23070 = x_reg_L0_31__retimed_I13052_QOUT;
reg x_reg_L0_31__retimed_I13049_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13049_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[12];
	end
assign N23060 = x_reg_L0_31__retimed_I13049_QOUT;
reg x_reg_L0_31__retimed_I13046_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13046_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[11];
	end
assign N23050 = x_reg_L0_31__retimed_I13046_QOUT;
reg x_reg_L0_31__retimed_I13041_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13041_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[8];
	end
assign N23035 = x_reg_L0_31__retimed_I13041_QOUT;
reg x_reg_L0_31__retimed_I13035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13035_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[5];
	end
assign N23018 = x_reg_L0_31__retimed_I13035_QOUT;
reg x_reg_L0_31__retimed_I13032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13032_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[10];
	end
assign N23008 = x_reg_L0_31__retimed_I13032_QOUT;
reg x_reg_L0_31__retimed_I13025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13025_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[4];
	end
assign N22989 = x_reg_L0_31__retimed_I13025_QOUT;
reg x_reg_L0_31__retimed_I13022_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13022_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[1];
	end
assign N22979 = x_reg_L0_31__retimed_I13022_QOUT;
reg x_reg_L0_31__retimed_I13019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13019_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[2];
	end
assign N22969 = x_reg_L0_31__retimed_I13019_QOUT;
reg x_reg_L0_31__retimed_I13016_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13016_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[3];
	end
assign N22959 = x_reg_L0_31__retimed_I13016_QOUT;
reg x_reg_L0_31__retimed_I13013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13013_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[9];
	end
assign N22949 = x_reg_L0_31__retimed_I13013_QOUT;
reg x_reg_L0_31__retimed_I13010_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13010_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[7];
	end
assign N22939 = x_reg_L0_31__retimed_I13010_QOUT;
reg x_reg_L0_31__retimed_I13007_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I13007_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[6];
	end
assign N22929 = x_reg_L0_31__retimed_I13007_QOUT;
reg x_reg_L0_31__retimed_I12919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12919_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365;
	end
assign N22618 = x_reg_L0_31__retimed_I12919_QOUT;
reg x_reg_L0_31__retimed_I12818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12818_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102;
	end
assign N22309 = x_reg_L0_31__retimed_I12818_QOUT;
reg x_reg_L0_31__retimed_I12816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12816_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240;
	end
assign N22305 = x_reg_L0_31__retimed_I12816_QOUT;
reg x_reg_L0_31__retimed_I12715_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12715_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944;
	end
assign N22003 = x_reg_L0_31__retimed_I12715_QOUT;
reg x_reg_L0_31__retimed_I12713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12713_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075;
	end
assign N21999 = x_reg_L0_31__retimed_I12713_QOUT;
reg x_reg_L0_31__retimed_I12711_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12711_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437;
	end
assign N21993 = x_reg_L0_31__retimed_I12711_QOUT;
reg x_reg_L0_31__retimed_I12710_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12710_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298;
	end
assign N21988 = x_reg_L0_31__retimed_I12710_QOUT;
reg x_reg_L0_31__retimed_I12644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12644_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246;
	end
assign N21795 = x_reg_L0_31__retimed_I12644_QOUT;
reg x_reg_L0_31__retimed_I12639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12639_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328;
	end
assign N21782 = x_reg_L0_31__retimed_I12639_QOUT;
reg x_reg_L0_31__retimed_I12634_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12634_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055;
	end
assign N21769 = x_reg_L0_31__retimed_I12634_QOUT;
reg x_reg_L0_31__retimed_I12632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12632_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188;
	end
assign N21765 = x_reg_L0_31__retimed_I12632_QOUT;
reg x_reg_L0_31__retimed_I12380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12380_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950;
	end
assign N21105 = x_reg_L0_31__retimed_I12380_QOUT;
reg x_reg_L0_31__retimed_I12378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12378_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362;
	end
assign N21100 = x_reg_L0_31__retimed_I12378_QOUT;
reg x_reg_L0_31__retimed_I12374_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12374_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115;
	end
assign N21090 = x_reg_L0_31__retimed_I12374_QOUT;
reg x_reg_L0_31__retimed_I12372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12372_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927;
	end
assign N21085 = x_reg_L0_31__retimed_I12372_QOUT;
reg x_reg_L0_31__retimed_I12370_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12370_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335;
	end
assign N21080 = x_reg_L0_31__retimed_I12370_QOUT;
reg x_reg_L0_31__retimed_I12368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12368_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901;
	end
assign N21075 = x_reg_L0_31__retimed_I12368_QOUT;
reg x_reg_L0_31__retimed_I12366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12366_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138;
	end
assign N21070 = x_reg_L0_31__retimed_I12366_QOUT;
reg x_reg_L0_31__retimed_I12237_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12237_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976;
	end
assign N20660 = x_reg_L0_31__retimed_I12237_QOUT;
reg x_reg_L0_31__retimed_I12190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12190_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400;
	end
assign N20538 = x_reg_L0_31__retimed_I12190_QOUT;
reg x_reg_L0_31__retimed_I12181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12181_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22];
	end
assign N20492 = x_reg_L0_31__retimed_I12181_QOUT;
reg x_reg_L0_31__retimed_I12116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12116_QOUT <= a_exp[5];
	end
assign N20182 = x_reg_L0_31__retimed_I12116_QOUT;
reg x_reg_L0_31__retimed_I12113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12113_QOUT <= a_exp[6];
	end
assign N20175 = x_reg_L0_31__retimed_I12113_QOUT;
reg x_reg_L0_31__retimed_I12103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12103_QOUT <= a_exp[0];
	end
assign N20144 = x_reg_L0_31__retimed_I12103_QOUT;
reg x_reg_L0_31__retimed_I12021_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12021_QOUT <= a_exp[1];
	end
assign N19909 = x_reg_L0_31__retimed_I12021_QOUT;
reg x_reg_L0_31__retimed_I12017_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12017_QOUT <= a_exp[2];
	end
assign N19900 = x_reg_L0_31__retimed_I12017_QOUT;
reg x_reg_L0_31__retimed_I12013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I12013_QOUT <= a_exp[4];
	end
assign N19891 = x_reg_L0_31__retimed_I12013_QOUT;
reg x_reg_L0_31__retimed_I11972_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11972_QOUT <= a_exp[3];
	end
assign N19768 = x_reg_L0_31__retimed_I11972_QOUT;
reg x_reg_L0_31__retimed_I11920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11920_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647;
	end
assign N19633 = x_reg_L0_31__retimed_I11920_QOUT;
reg x_reg_L0_31__retimed_I11828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11828_QOUT <= a_man[0];
	end
assign N19410 = x_reg_L0_31__retimed_I11828_QOUT;
reg x_reg_L0_31__retimed_I11770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11770_QOUT <= a_man[1];
	end
assign N19275 = x_reg_L0_31__retimed_I11770_QOUT;
reg x_reg_L0_31__retimed_I11753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11753_QOUT <= a_man[3];
	end
assign N19233 = x_reg_L0_31__retimed_I11753_QOUT;
reg x_reg_L0_31__retimed_I11749_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11749_QOUT <= a_man[2];
	end
assign N19223 = x_reg_L0_31__retimed_I11749_QOUT;
reg x_reg_L0_31__retimed_I11721_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11721_QOUT <= a_man[7];
	end
assign N19159 = x_reg_L0_31__retimed_I11721_QOUT;
reg x_reg_L0_31__retimed_I11717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11717_QOUT <= a_man[10];
	end
assign N19149 = x_reg_L0_31__retimed_I11717_QOUT;
reg x_reg_L0_31__retimed_I11713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11713_QOUT <= a_man[6];
	end
assign N19139 = x_reg_L0_31__retimed_I11713_QOUT;
reg x_reg_L0_31__retimed_I11709_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11709_QOUT <= a_man[8];
	end
assign N19129 = x_reg_L0_31__retimed_I11709_QOUT;
reg x_reg_L0_31__retimed_I11705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11705_QOUT <= a_man[11];
	end
assign N19119 = x_reg_L0_31__retimed_I11705_QOUT;
reg x_reg_L0_31__retimed_I11701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11701_QOUT <= a_man[12];
	end
assign N19109 = x_reg_L0_31__retimed_I11701_QOUT;
reg x_reg_L0_31__retimed_I11697_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11697_QOUT <= a_man[13];
	end
assign N19099 = x_reg_L0_31__retimed_I11697_QOUT;
reg x_reg_L0_31__retimed_I11689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11689_QOUT <= N30313;
	end
assign N19080 = x_reg_L0_31__retimed_I11689_QOUT;
reg x_reg_L0_31__retimed_I11685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11685_QOUT <= a_man[5];
	end
assign N19070 = x_reg_L0_31__retimed_I11685_QOUT;
reg x_reg_L0_31__retimed_I11681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11681_QOUT <= a_man[9];
	end
assign N19060 = x_reg_L0_31__retimed_I11681_QOUT;
reg x_reg_L0_31__retimed_I11677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11677_QOUT <= a_man[14];
	end
assign N19050 = x_reg_L0_31__retimed_I11677_QOUT;
reg x_reg_L0_31__retimed_I11673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11673_QOUT <= a_man[15];
	end
assign N19040 = x_reg_L0_31__retimed_I11673_QOUT;
reg x_reg_L0_31__retimed_I11669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11669_QOUT <= a_man[18];
	end
assign N19030 = x_reg_L0_31__retimed_I11669_QOUT;
reg x_reg_L0_31__retimed_I11665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11665_QOUT <= a_man[20];
	end
assign N19020 = x_reg_L0_31__retimed_I11665_QOUT;
reg x_reg_L0_31__retimed_I11661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11661_QOUT <= a_man[17];
	end
assign N19010 = x_reg_L0_31__retimed_I11661_QOUT;
reg x_reg_L0_31__retimed_I11657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11657_QOUT <= a_man[19];
	end
assign N19000 = x_reg_L0_31__retimed_I11657_QOUT;
reg x_reg_L0_31__retimed_I11653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11653_QOUT <= a_man[16];
	end
assign N18990 = x_reg_L0_31__retimed_I11653_QOUT;
reg x_reg_L0_31__retimed_I11645_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11645_QOUT <= a_man[21];
	end
assign N18971 = x_reg_L0_31__retimed_I11645_QOUT;
reg x_reg_L0_22__retimed_I11608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I11608_QOUT <= a_man[22];
	end
assign N18886 = x_reg_L0_22__retimed_I11608_QOUT;
reg x_reg_L0_31__retimed_I11606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11606_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577;
	end
assign N18881 = x_reg_L0_31__retimed_I11606_QOUT;
reg x_reg_L0_31__retimed_I11605_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11605_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487;
	end
assign N18879 = x_reg_L0_31__retimed_I11605_QOUT;
reg x_reg_L0_23__retimed_I11588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I11588_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580;
	end
assign N18839 = x_reg_L0_23__retimed_I11588_QOUT;
reg x_reg_L0_23__retimed_I11586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I11586_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026;
	end
assign N18835 = x_reg_L0_23__retimed_I11586_QOUT;
reg x_reg_L0_16__retimed_I11519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I11519_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82;
	end
assign N18678 = x_reg_L0_16__retimed_I11519_QOUT;
assign N30269 = !N18678;
assign N30270 = !N30269;
reg x_reg_L0_21__retimed_I11514_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I11514_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759;
	end
assign N18667 = x_reg_L0_21__retimed_I11514_QOUT;
assign N30271 = !N18667;
assign N30276 = !N30271;
assign N30275 = !N30271;
assign N30274 = !N30271;
assign N30273 = !N30271;
assign N30272 = !N30271;
reg x_reg_L0_31__retimed_I11513_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11513_QOUT <= a_sign;
	end
assign N18664 = x_reg_L0_31__retimed_I11513_QOUT;
reg x_reg_L0_31__retimed_I11511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I11511_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639;
	end
assign N18660 = x_reg_L0_31__retimed_I11511_QOUT;
assign N30277 = !N18660;
assign N30284 = !N30277;
assign N30283 = !N30277;
assign N30282 = !N30277;
assign N30281 = !N30277;
assign N30280 = !N30277;
assign N30279 = !N30277;
assign N30278 = !N30277;
assign bdw_enable = !astall;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316 = ((a_exp[4] & a_exp[3]) & a_exp[5]) & a_exp[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639 = !(a_exp[7] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13316);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360 = !a_exp[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345 = !a_exp[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349 = !(a_exp[2] & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347 = !(a_exp[4] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5347) ^ a_exp[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5349) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5360;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1] = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5345;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1] ^ a_exp[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0] = !a_exp[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595 = !a_man[21];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595 | a_man[19];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168} = {1'B0, a_man[17]} + {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4489};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181 = !a_man[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181 | a_man[20];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374} = {1'B0, a_man[18]} + {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4153} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4212} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4374};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181) ^ a_man[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274 = !a_man[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274 | a_man[18];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064} = {1'B0, a_man[16]} + {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4113};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4554} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3994} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4168};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595) ^ a_man[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958 = !a_man[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958 | a_man[17];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959} = {1'B0, a_man[15]} + {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4449};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4176} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4331} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4064};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274) ^ a_man[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368 = !a_man[18];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368} + {1'B0, a_man[13]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577} = {1'B0, a_man[14]} + {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4387};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4516} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3953} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3959};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958) ^ a_man[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052 = !a_man[17];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166} = {1'B0, a_man[12]} + {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571} = {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4319} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4012};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4141} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4294} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4577};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454 = !a_man[16];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4571} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3943} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4166};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4075} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4229} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4471};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548 = !a_man[14];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403} = {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145 = !a_man[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342} = {1'B0, a_man[22]} + {1'B0, a_man[13]} + {1'B0, a_man[10]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4215} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4560} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4342};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989} = {1'B0, a_man[11]} + {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4283};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4438} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4378} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4109};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4504} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4411} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4600};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360} = {1'B0, a_man[12]} + {1'B0, a_man[9]} + {1'B0, a_man[7]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144} = {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608} = {1'B0, a_man[8]} + {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4297};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4493} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4403} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4360};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4307} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4156};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4348} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3989};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236 = !a_man[13];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271} = {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014} = {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118} = {1'B0, a_man[7]} + {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4169};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4366} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4592} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4608};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4427} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4026} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4334};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4061} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4224};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922 = !a_man[12];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613} = {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958};
assign N30312 = !a_man[4];
assign N30313 = !N30312;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351} = {1'B0, a_man[6]} + {1'B0, N30313} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4041};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4235} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4453} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4118};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4271} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4623} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4204};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4247} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4001} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4243};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322 = !a_man[11];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596} = {1'B0, a_man[5]} + {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4613};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4103} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4321} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4351};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4144} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4483} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4076};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4120} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4180} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4478};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015 = !a_man[10];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220} = {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4193} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4219} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4596};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4014} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4352} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3946};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3985} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4050} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3999};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457} = {1'B0, a_man[6]} + {1'B0, a_man[3]} + {1'B0, a_man[1]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104 = !a_man[8];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584} = {1'B0, a_man[22]} + {1'B0, a_man[15]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4249} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4006} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4220};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415 = !a_man[9];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415} + {1'B0, N30313};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4183} + {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4106};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3970} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4065} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4532};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4574} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3919} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4232};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508 = !a_man[7];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4029} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4369} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4584};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456} = {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604} = {1'B0, a_man[5]} + {1'B0, a_man[2]} + {1'B0, a_man[0]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4121} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4624} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4457};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4564} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4090} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4636};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4507} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4440} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4468};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080 = !a_man[6];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923} = {1'B0, a_man[13]} + {1'B0, N30313} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4170} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4079} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3995};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4456} + {1'B0, a_man[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4604};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3960} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4207} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4404};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4469} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4380} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3987};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614 = !a_man[5];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230} = {1'B0, a_man[1]} + {1'B0, a_man[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4355};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4549} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4524} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4053};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4597} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3935} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4338};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158} = {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494} = {1'B0, a_man[3]} + {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4638};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4107} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4016} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4230};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4289} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4194} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4494};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4441} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3923} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3948};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4300} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4392} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4476};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428 = !a_man[3];
assign N30285 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428;
assign N30286 = !N30285;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104} + {1'B0, N30286};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4032} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3938} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4158};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287 = !a_man[4];
assign N30287 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287;
assign N30288 = !N30287;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039} = {1'B0, a_man[11]} + {1'B0, N30288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069} = {1'B0, a_man[2]} + {1'B0, a_man[17]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4039};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4383} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4472} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4221};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4238} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4580} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4115};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056} = {1'B0, a_man[9]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393} = {1'B0, a_man[1]} + {1'B0, a_man[16]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4210};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4406} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4314} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4069};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4510} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4134} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4377};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381 = !a_man[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488 = a_man[15] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4488};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3963} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4601} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4393};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4149} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4056} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3936};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4303} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4499} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4526};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4162} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4251} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3920};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316 = (!a_man[15]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4197} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4267} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4316};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198} = {1'B0, a_man[8]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417 = !a_man[1];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4198};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4241} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4329} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4083};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4093} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4432} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4276};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227} = {1'B0, a_man[13]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4181};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4139} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4386} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4557};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084} = {1'B0, a_man[14]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4112} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4174};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3992} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4371} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4533};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949 = !a_man[0];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336} = {1'B0, a_man[5]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4099} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4318} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4227};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4047} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3976};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4020} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4084};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410} = {1'B0, a_man[12]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575} = {1'B0, N30313} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4410} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4502} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4336};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983} = {1'B0, N30288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4569} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4165};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3952} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4619} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4437};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607} = {1'B0, a_man[11]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4274};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092} = {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4607} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3967} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4575};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218} = {1'B0, N30286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4035} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4347};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4073} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4539} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3983};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059} = {1'B0, a_man[10]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3958};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326} = {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4059} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4155} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4092};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4213} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4529};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4254} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4010} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4218};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4621);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087 = a_man[9] | N30288;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931 = (!a_man[9]) ^ N30288;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3931};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4087} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4632};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4189} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4436} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4455};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343} = {1'B0, a_man[8]} + {1'B0, N30286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4052};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4024} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4490} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4326};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4376} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3997} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3971};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3984);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049} = {1'B0, a_man[7]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4454} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4519} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4202} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4343};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4591} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4556} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4208};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4463;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4128;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481 = a_man[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4481};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982} = {1'B0, a_man[6]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4145};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4049} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4143};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4622} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4365} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4461};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4270} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4425} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4225};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4548} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3982} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4543} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4587};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609} = {1'B0, N30313} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4236} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320 = (!a_man[5]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4320} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4167} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3978};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119} = {1'B0, a_man[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4322};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998} = {1'B0, a_man[3]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3945} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3998};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4412} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4609};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350} = {1'B0, a_man[0]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4415};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233} = {1'B0, a_man[1]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4015} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4439} + {1'B0, N30288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4233};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4191} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4119};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4104} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4379} + {1'B0, N30286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4350};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4508} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4080};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4467} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4217};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635} = {1'B0, N30288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4308};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004} = {1'B0, N30286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949} + {1'B0, a_man[6]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4614} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4287} + {1'B0, N30286};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4428;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961 = !(a_man[1] | a_man[0]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4381;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3949 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4273);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4071 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4385) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4226);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3961) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4184)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4030);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4417 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4182);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4496 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4335);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4537 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4137;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3975) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4312) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4617) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4578)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3933) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4004));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4157 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4635);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4205 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4196) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4045);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4513) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4563)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4063) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3968 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4131);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4284 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4611);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3951 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4265;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4420 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4110) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4101) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4546);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4559) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4491);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4038 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4349);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4505 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4100);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4582 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4327) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4173);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4257 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4573);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4013 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4231);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4486 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4239) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4081);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4401) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4464)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4306);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4266 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4583;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4389 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4296);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4450 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3955);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4396 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3990;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4148 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4550) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4330) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3944);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4117 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4177);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4333 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4305);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4301 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4054) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4443) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4512)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4356);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19007) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3918)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19009) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19011));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4281 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3941);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4542 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4295) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4097 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4477)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4111) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4585)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4422);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4641 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4292);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4451 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4203) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4446 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4421)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4586 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4397);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4552 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4124)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4487)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4328);
assign N30315 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4008;
assign N30316 = (!N30315) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4161 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042 = !N30316;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4278 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4567);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4007 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4535)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3972 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4263);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4416 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3988)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4398)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4240);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4146 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4275);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4430 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4160)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4309 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4132);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4285 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4259)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4302)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4150);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4068) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4637);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4509)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4354);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4413 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4390);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4521)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3957 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3932);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4088 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4465)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4209)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4055);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4634 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4610);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4036 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4098)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4256 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4479);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4540 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3917)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4125)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3962);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4534;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3973 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4324);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3979 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4201);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4361 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4588)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4022 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4400 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4630)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4031)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4602);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4206)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4280 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4200)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4363);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025} = {1'B0, a_man[22]} + {1'B0, a_man[19]} + {1'B0, a_man[17]};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4528} + {1'B0, a_man[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4025};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4515) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4424 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344} = {1'B0, a_man[20]} + {1'B0, a_man[18]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4187};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4228);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4538) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4434 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4605)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4523 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4102) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4258);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4344 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4034);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4423)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4590);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940} = {1'B0, a_man[21]} + {1'B0, a_man[19]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4021) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4414 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4255;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4480)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4074) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4011;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4268 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4409;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4431;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4277;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4199 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4612) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4040);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4164;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3981)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4140);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4293) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4640;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4192 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4317;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152 = (!a_man[22]) ^ a_man[21];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253} = {1'B0, a_man[22]} + {1'B0, a_man[20]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4138);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4339);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4288);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3977 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4447) | (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3940 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4501)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4185) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3937)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4498);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4133 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4615) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4484) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4418)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4262);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4095 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4253);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4595 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4408) & (!(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359)));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4482);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152) & (a_man[22] | a_man[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4122;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4618;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3929)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4085);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4244) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4359;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4589 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4046;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3921) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4152;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5348 ^ a_exp[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5489);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5478 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5415 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5506 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign N30323 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5524);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778 = !N30323;
assign N30289 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778;
assign N30293 = !N30289;
assign N30292 = !N30289;
assign N30291 = !N30289;
assign N30290 = !N30289;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N750) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N631 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N630 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N633 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N632 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N627 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N626 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N629 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N628 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N635 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N637 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N636 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5389);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N751) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5443 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5534 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5451 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5425 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5500);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N752) ^ N30293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5460 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5553 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5486 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5581 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5434);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5400);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N753) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5778;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5544 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5570 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5397 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5513);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N754) ^ N30293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5377 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5404 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5413);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N755) ^ N30293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6006 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5891);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[20];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6076 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6130 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6456);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[22]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[17] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6187 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6299 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6008);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5957 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6633 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6171) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5869) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6057);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5868);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6087);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5988);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6248) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6355) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6521);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6317 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6667;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6004;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6614);
assign N30329 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180 = !N30329;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6127) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6018) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6197 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6552) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6483));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255 = 1'B0 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6574 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6300);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5885 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6365 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6440;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5974;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6002 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6264);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6538) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6618) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5890);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[27] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6156 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6509) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6074));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[27]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6466 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5923;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5905;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6106 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6141) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5959) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6391);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[26] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5927 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6033) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[26]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391 = N29673 & N29667;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6215 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6605;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5907;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6635;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6458;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6555;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6568 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6437;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6366;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6389;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6022;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6201 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6557) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6285) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6095);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[25] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6174 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6357) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6525) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5994);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929} = {1'B0, 1'B1} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[25]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4382) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4222);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4525)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4372);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4346);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4570 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4096;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3969) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4503;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5561 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5530 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5548 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5477);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N748) ^ N30293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4299;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3942 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4188;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N625 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N624 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5432 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5483 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5501 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N747) ^ N30293;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5516 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5395 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5525 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5497 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5378);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N749 ^ N30292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8982;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42] = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9472 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5840 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6540 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6159 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6442);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5861 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6237) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6407) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5945);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042);
assign N30373 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6511;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 = !N30373;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6591 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6131));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8770) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6380;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6284;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5944;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6513;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6185;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6172;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6496;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5980 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37720);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6408;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6670;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6217;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6266;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6422;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6343;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6160) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6347) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5862);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[24] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6132 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6318) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6485) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5946);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[24]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[41] = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[42];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6195;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6663;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5902;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6473 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6301) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6654) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6009;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[23] = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6077 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6189) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6543) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6368;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5522);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4114) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4606;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N622 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5468 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5385 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5455 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5454);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N746) ^ N30292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4579;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4628)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4459);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4530);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4037 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4282;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5422 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5552 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5392 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5433 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5408 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5407);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N745) ^ N30292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9016;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9506 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8794) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6542 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6443) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6078) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6270);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8822) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[41], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[40]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9163};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[23]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[41]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[41]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6334;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5846;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6499;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6154;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6481;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6550;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6258 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5965) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6609) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6145);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[22] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6221 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6395) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6577) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6036);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5842;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6396 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5931) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6576);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8881) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9700;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8849) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5550);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4066) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3966;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N620 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5375 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5504 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5558 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5505 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5575 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N744) ^ N30292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5457);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4048;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4631);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4129 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4375;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N619 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5542 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5459 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5511 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5579 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5529 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5528);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N743) ^ N30292;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9052;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6042) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6610) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6066) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5878);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6257 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5964));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8941) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9200} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10137};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[40], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[39]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9307} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8802} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9919};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12365} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[22]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[40]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[40]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11918 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12437;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391 & N29566;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6099;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6280;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6677) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6639) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5912);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[21] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5997 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6361) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6288));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9539 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8818) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3954) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4060;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N618 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5495 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5414 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5465 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5442 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5481 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5480);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N742) ^ N30291;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5576);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3991;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4473;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4313;
assign N30336 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4078)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4237));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394 = !N30336;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4551;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4565) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4005);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3996;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4633)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4062);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4214) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4462;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N617 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5449 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5578 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5420 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5437 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5436);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N741) ^ N30291;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9083;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8912) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9627} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8836};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8972) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8877) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9238} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10171} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9235};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6233;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6414) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6322) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6595);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6678) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5951) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6135);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9005) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9763} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9779} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9056} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8994};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[39], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[38]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9373} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9538} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10126};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12222, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12080} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[39]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[39]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970 = !(N22618 & N29506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5986;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6350;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6166;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6083) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6447) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6277);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[20] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6051 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6242) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6413) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5865);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9569 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8846) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4159 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4154;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N616 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5402 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5427 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5374 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5390 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5388);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N740) ^ N30291;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4394;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4086;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4402)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4562);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4000) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4558;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N615 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5567 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5485 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5381 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5539 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5448 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5556 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N739) ^ N30291;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9121;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8939) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9667} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8867};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6332;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6403) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6117);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6453;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6523;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6093;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6305) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6477) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5898) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6448)) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6012) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6084);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9067) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8844, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9392} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8769} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8718};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5970) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6149) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6339);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6406;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6502) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5851 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6227));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9128) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9033) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9002) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8910) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9271} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10206} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9299};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9814} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9010} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8694};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6089;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6492;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6387) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5838;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5918) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6028 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6212) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6566 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6102) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9194) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9095) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9600 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8875) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4517 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4246;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N614 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5521 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5441 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5547 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5492 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5509 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5508);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N738) ^ N30291;
assign N30343 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4082)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3928));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934 = !N30343;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4492 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3930;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N613 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5474 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5499 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5446 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5566 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5463 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5462);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N737) ^ N30290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9157;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8969) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9702} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8904};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9429} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8679} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10280};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9890} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10103} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10159} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9116};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9601, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9212} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9509} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10185} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10249};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[38], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[37]} = {1'B0, N23333} + {1'B0, N23335} + {1'B0, N29612};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446} = {1'B0, N23140} + {1'B0, N23142} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[38]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323 = !(N29502 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6630;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6451;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6340;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6310) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6616) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6306) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6478) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6228);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[19] = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6400 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5936) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6116) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6658;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9158) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9065) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6352 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6402) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6193) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6016;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6373;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6169) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5901 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6548) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6247 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5990) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6353) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6418);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9259) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9853} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9044} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9991};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9181, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8821} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9318} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10011} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9796};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6153) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6505) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6342);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5853 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6587) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6043) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6232);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9327) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9463} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8708} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9618};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9031) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8937) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9313} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10244} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9365};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10073, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8726} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10194} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9926};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9091) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8999) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9190) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8936} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9885} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9075};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9634 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8906) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3934) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4332;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N612 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5429 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5560 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5373 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5453 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5399 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5520 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5418 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5417);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N736) ^ N30290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4042;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4269);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4594 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4023;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N611 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5514 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5541 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5406 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5565 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5473 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5584 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N735) ^ N30290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9196;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5922) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6107) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6468);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6293 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6647) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6184) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6003);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6536 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5887;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9394) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9740} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9230};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8852} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8828} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9582} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10045};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9089, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8744} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8940} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9221} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9709};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574} = {1'B0, N23943} + {1'B0, N23945} + {1'B0, N29496};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909} = {1'B0, N23579} + {1'B0, N29498} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9954};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__115__W1[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[13];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7554} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7522} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7670};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7986};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7568} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7540} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7754};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8043} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7685} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7861};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7888} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7821} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7626};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[9];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7957} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8002} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7744};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7546} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7527} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7667};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7794} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7910} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8039};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7648} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7703} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7894};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[7];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8077} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7867} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8060};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7847} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8035} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7981};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7613} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7615} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7864};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7521} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7723} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7771};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7599} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7732} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7741};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7765} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8062} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7747};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7915} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7594};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8049} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7745} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7539};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7677} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7801} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8073};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7859} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8061} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7693};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8057} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7556} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7803};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7905} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7641} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7586};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7938} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7920} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7811};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7788} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7933} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7662};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8009} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7695} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7987};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7551} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7822} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7588};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7560} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7994} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7565};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7772} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8019} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8001};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7533} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7782} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8052};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7887} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7832} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7567};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7873} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7577} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7992};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7611} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7813} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7989};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7932} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7566} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7906};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7674} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7650} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7896};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7684} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7705} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7947};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8030} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7736} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7715};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4362) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4426;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N610 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5456 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5467 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5494 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5573 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5519 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5428 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5537 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5536);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N734) ^ N30290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1];
assign N30294 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958;
assign N30302 = !N30294;
assign N30301 = !N30294;
assign N30300 = !N30294;
assign N30299 = !N30294;
assign N30298 = !N30294;
assign N30297 = !N30294;
assign N30296 = !N30294;
assign N30295 = !N30294;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885 = N30302 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8068} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7624} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7885};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2];
assign N30303 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696;
assign N30311 = !N30303;
assign N30310 = !N30303;
assign N30309 = !N30303;
assign N30308 = !N30303;
assign N30307 = !N30303;
assign N30306 = !N30303;
assign N30305 = !N30303;
assign N30304 = !N30303;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007 = N30311 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7690} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7886} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7664};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8007} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7959} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7889};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582 = !(N30311 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7895} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7749} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7582};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7642} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7865} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7544};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7916} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7579} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7596};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7926} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7628} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7605};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7834} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8088} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7767};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7943} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7649} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7639};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059 = !(N30302 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4518;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4175;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4019;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4405 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4429) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4364;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4028) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4367)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N3956) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N4116;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N609 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[0]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N608 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5493));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5410 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5540) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5502 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5421 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5562) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5447 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5568));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5527 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5545) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5472 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5379));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5382 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[4]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5488);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N733 ^ N30290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900 = !(N30311 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7977} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7764} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7900};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7687} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7606} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7855};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7569} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7815} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7793};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7824} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7843} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8075};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8059) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8065;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7724} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7702};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7967} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7737};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7652} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7558} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7580};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809 = !(N30302 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655 = !(N30311 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7762} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7809} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7655};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7898} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8054} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7738};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7534} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8011} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7783};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8041} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8064} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7727};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564 = !(N30301 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7564} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7570};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7955} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7868} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7524};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7875);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7770} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7791};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7714} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8053} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7515};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8000);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971 = !(N30311 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7725} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8038} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7971};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7548} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7796} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8021};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7826} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7978} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8078};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7697} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8031} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7936};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730 = !(N30310 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8040} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7890} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7730};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884 = !(N30301 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7884} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8029} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7804};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7750} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7768} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8013};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7774} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8044} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7706};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7665} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7757} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7907};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637 = !(N30301 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7637} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7643};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7755);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7542} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7557};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7983} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7962} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7668};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7993} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7675} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7698};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7729} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7949} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7631};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7627);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7862} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7543};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046 = !(N30310 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8046} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7881} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7858};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7644} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7912} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7891};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7918} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7939} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7598};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713 = !(N30301 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7713} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7718};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7532} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7877} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8024};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954 = !(N30301 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798 = !(N30310 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7961} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7954} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7798};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7561} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7806} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7537};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7571} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7591} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7817};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7575);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8074);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549 = !(N30310 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7616} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7630} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7549};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7760} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7710} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8005};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7786} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8058} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8034};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7946);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7935} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7617};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027 = !(N30300 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8033} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8027} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7948};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7601} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7901} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7848};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7689} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7930};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7958 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7780} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7785};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870 = !(N30310 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7870} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7996} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8047};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7528} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7583} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7828};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621 = !(N30309 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7823);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8010} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7536};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7694} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7621} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7819};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7731} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7972};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531 = !(N30300 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941 = !(N30309 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7531} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8020} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7941};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7871} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8069} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7550};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851 = !(N30300 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7578);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7851} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7766};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7892} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7700} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7942};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7842);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8084} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7608};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699 = !(N30309 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7699} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7965} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7769};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014 = !(N30309 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604 = !(N30300 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7604} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8014} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7840};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925 = !(N30300 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7726);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7925} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7833};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7990);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681 = !(N30299 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7696);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7587} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7681};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517 = !N30309;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | N30299) | N30308);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7850) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7612)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7914));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8037 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7593);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7721 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7530) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7974);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7779) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7573)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7722) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7518));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7646 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8015);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7921 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8026) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7903);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7712) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7709)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7574) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7622));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7752 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7799);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7922 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7656);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7830 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8083);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7911;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7636 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7953) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7982) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7520);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7883) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7795)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7777) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8081));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7634 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7609);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7742 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7719);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8006 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7692;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7808 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7686) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19018 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7673) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7838 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8066);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7619 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7844);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7970 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7878);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8016 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7820) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7701);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7931) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7743)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7610);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8003 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7589);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7716 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7618);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7623);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7748 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7968);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7523 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7756);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7552);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7669)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7538);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7940) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7818);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7876 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7853);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7976 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7956);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8048);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8086 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7814);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7934 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7672);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7973);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7592)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8036);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7790 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7841);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7966 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8017);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7902);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7945 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7576);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8072 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7874);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7829);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7516)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7963);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7869) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7751);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7797)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7553 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7998);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7802 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7680);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7761);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7645;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7929);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7789) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7924));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7555 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7683));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[32] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8076) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7807;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[31] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8056) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7825;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468} = {1'B0, N29614} + {1'B0, N29598};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10214;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9468;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[37], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[36]} = {1'B0, N29610} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9279} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10192};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164} = {1'B0, N23130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[37]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[37]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37712);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6133;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6182;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5917) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6292) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6103);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[18] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5882 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6261) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6534);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5942 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6125) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6313) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6664);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8851 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6482 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6017));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692 = ((!N30268) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9061) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8964) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9347} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10276} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9433};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9289) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6522) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5870) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6058);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6140) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6250) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6603) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6420);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9459) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9155) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9256) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9503} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8859} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8738};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10027} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9162} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8945};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9668 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[3]) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8934) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9424) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134} = {1'B0, N30308} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9774} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9266};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9357) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9122) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9028) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9222) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8971} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9923} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9111};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9660} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9526} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10263};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10165} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9191} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9716};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9983, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9611} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9835} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8648} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9354};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9325) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6128 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6315) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6484) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6668);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6554) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6020) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6378) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6199);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9528) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9088) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8997) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9386} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10307} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7517};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10199} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10059} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10089};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8801} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10286} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9294};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10109, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9746} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9960} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8748} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8977};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671} = {1'B0, N24432} + {1'B0, N29490} + {1'B0, N29655};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478} = {1'B0, N29492} + {1'B0, N29494} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9004};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6073 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6267) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6438) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6537);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10191 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6155) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6617) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5975);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925 = ((!N30266) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30268));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9574} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9862} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8925};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[36], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[35]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8909} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9692} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8967};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522} = {1'B0, N23120} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[36]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[36]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7846;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8082;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7651)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7773);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[30] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7897) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7882;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[29] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7810 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7635;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596 = !(N29592 | N29580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9596 | N29598;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6032 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6218) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6570) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6497);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9832 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6109) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5924) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6390);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909 = ((!N30264) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6075) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6269) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6619);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5978) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5858) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6441) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6345) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6157);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9592) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9390) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[1] & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993 | (!N30299));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8962) & N30308));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9693} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9844} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9913};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9187) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9286) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9541} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8896} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8762};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9687} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9877} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8895} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9134};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9486, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9098} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10050} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9326} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10079};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9559) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026 = !((N30299 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664) | ((!N30299) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9026) & N30308));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9766} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9421};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9355) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9732} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10235} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10098};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9152) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9058) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9253) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9007} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9955} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9148};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9265} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9695} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8737} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9726};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9072, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8731} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9904} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9659} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8919};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9808) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9302;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6034) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5843) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5928);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6219) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6298) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6392) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6573);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9662) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9218) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9119) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8673} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9576} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9340};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9457} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9530} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8764};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8710, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10026} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9496} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10234} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9462};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456} = {1'B0, N25766} + {1'B0, N25768} + {1'B0, N29486};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869} = {1'B0, N29488} + {1'B0, N29624} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9843};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776} = {1'B0, N29626} + {1'B0, N29653} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10229};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9447 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5872 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6423) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6251);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137 = ((!N30262) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30264));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8671} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9127} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9137};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9478} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9909} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9771};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[35], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[34]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10303} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8880};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6417 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6599) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6325) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5953);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[17] = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6493 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6137));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245} = {1'B0, N23110} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[35]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[35]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6374 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6549) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5900) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6088;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[16] = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5991 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6452) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6060;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251 = (!N29598) | (N29592 & N29580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10251;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 = (!N29592) ^ N29580;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8992) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7839;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7620;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8067;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7919)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8045);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7720;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7633) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7759);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7584;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8042)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[28] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7728) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7952;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[27] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7880 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7711;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495 = !(N29426 | N29570);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9495 | N29580;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5855 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5888) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6671) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6094) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9064 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6556 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6457;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118 = ((!N30260) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9525) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5908;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5995;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6200 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6547) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6649) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5874) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6062) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6636);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6175 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6359) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6527) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6254);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9728) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9322) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9070} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8793};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10208, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9852} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9502} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9301} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10058};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043} = {1'B0, N26244} + {1'B0, N26246} + {1'B0, N26248};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9387) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9690) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10267} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10129} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9493};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9184) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086 = !((N30299 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978) | ((!N30299) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8664));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9086) & N30308));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9283) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9040} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9986} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9186};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8903} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10278} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9312} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10097};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9624) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9420) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9847) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6409) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6239) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5947) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6592);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6672 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6486;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9788) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9376} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9338} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8732};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9733} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9878} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9540};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9237, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8866} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10243} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9274} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9078};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9756) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9250) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6079 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6544 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5893) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6272);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9854) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9613} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9102} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10051};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150 = !((N30298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599) | ((!N30298) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9150) & N30307));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9978);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8824;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8702} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10216};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9353) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9556) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9658) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8961} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8823} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9914};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9799} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9575} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10306};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10035, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9666} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9110} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10068} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9886};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629} = {1'B0, N26206} + {1'B0, N26208} + {1'B0, N29478};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816} = {1'B0, N29480} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9043} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9999};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9428} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9456} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10170};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7600;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7657;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7866)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7991);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[26] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7545) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8025;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[25] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7691 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7778;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396 = !(N29560 | N29430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9396 | N29570;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9869} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8858} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8776} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10118} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9257};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9382} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9896};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[34], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[33]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10067} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10221} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8796};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977} = {1'B0, N23100} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[34]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[34]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6615;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6044;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6265) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6436) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5973);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6504) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5886);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5941 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6123) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6588) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5854);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[15] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6231 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6311;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9114) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319 = (!N29580) | (N29426 & N29570);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9319;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 = (!N29426) ^ N29570;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8902) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9118} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9309} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9518};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[33], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[32]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9699} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10132} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8915};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329} = {1'B0, N23090} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[33]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[33]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6216 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6108) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6569) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6294;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign N30352 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648 = !N30352;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[14] = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5921 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6183) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6467) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6648;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6188) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6541);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6312 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6152) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6007;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6236 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6512) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5892) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5979) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5860);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363 = ((!N30258) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8959) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9363} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8887} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8768};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6428) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6608) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6144);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490);
assign N30360 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845 = !N30360;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10044 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6220) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5963) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6498) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5845);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659 = ((!N30256) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30258));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9085, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8742} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9149} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9922} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8935};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9418) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9621) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9724) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10300} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10161} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9531};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9739} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8672} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9414} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9185};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216 = !((N30298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208) | ((!N30298) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9216) & N30307));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9522) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8854;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9377} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10018} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10275};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9452) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9320) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9819) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6611 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6335) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5847) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6500);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6222) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6146) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6038);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9915) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8756} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9223} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9685};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9765} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9838} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9612};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9860, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9469} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9348} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10105} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9703};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714} = {1'B0, N26236} + {1'B0, N26238} + {1'B0, N29484};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9587) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9786) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9883) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9138} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8998} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10087};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9599);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281 = !((N30298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842) | ((!N30298) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9208));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9281) & N30307));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9297} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9654};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9384) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6562) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5913) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6460);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6178) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6289) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9976) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9688) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9295} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8855} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9948};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9872} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8890} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9653};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9120, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8771} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9956} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9385} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8970};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218} = {1'B0, N26198} + {1'B0, N29476} + {1'B0, N29482};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434} = {1'B0, N25627} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8873} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8714};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9051} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9629} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9823};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7913)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7787);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7733);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[24] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7937 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7529;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[23] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7708) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7849;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291 = !(N29442 | N27939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9291 | N29430;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9816} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9019} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8659} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10201} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9201};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9620} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8933} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9650};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[32], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[31]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10017} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10256} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9037};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054} = {1'B0, N23080} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[32]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[32]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6356 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5871) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6059) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[13] = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6331 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6249) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6421) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6604;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6206) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6382) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6560);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5911 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9677 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6638) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6098) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6287);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595 = ((!N30254) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110 = (!N29570) | (N29560 & N29430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10110;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 = (!N29560) ^ N29430;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8869) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9595} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8835} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9547};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6165) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6082 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N37704);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6276 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6274) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6446);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9284 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5950) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6241)) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6625) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5984);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839 = ((!N30244) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30254));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10134, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9773} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9450} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9224} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9985};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5987 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6031) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6449) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6517);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6628) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6243);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6053 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5952);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6167 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19032);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10036) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9655) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9754) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8667} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8920} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9568};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9039} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9689} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9489} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10231};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9554) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9907;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9413} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8666};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9484) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349 = !((N30298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183) | ((!N30298) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8842));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9349) & N30307));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9946) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8787} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9261} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9727};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10021} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9800} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9135} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8922};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9156, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8798} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8701} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9423} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9006};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511} = {1'B0, N26758} + {1'B0, N26760} + {1'B0, N29456};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9617) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9817) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9171;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9176} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9032} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8719};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9449) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9911) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10004) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9720) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9333} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10121} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9981};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10195} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10146} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9944};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6307 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6041) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6229) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5937);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6479) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6585) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6119);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10099) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415 = !((N30298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825) | ((!N30298) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9415) & N30307));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9519) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8888} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10261} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9836};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9073} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8955} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8783} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10264};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10167, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9807} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9260} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8733} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9460};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551} = {1'B0, N26654} + {1'B0, N29468} + {1'B0, N29454};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252} = {1'B0, N29474} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9511} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9928};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9891} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10218} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8911};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6040 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6226) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6399) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6582);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5969);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8914 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6304) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6114) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5935);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821 = ((!N30252) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30244));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9434} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9636} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9821};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8839} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8683} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8840};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9082) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9316) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9738} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9787} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9921};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9229} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9967} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8981};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9023) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8811) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9248) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9927} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10102} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10273};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[31], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[30]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9391} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8699};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416} = {1'B0, N23070} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[31]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[31]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161 = (!N29430) | (N29442 & N27939);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9161;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 = (!N29442) ^ N27939;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8734) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8929) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9146) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9154} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8976} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9345};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8810} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9591} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8656};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[30], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[29]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9990} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9753} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9012};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6129 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6669) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6316) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[12] = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6021 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6092) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6379) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6198;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132} = {1'B0, N23060} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[30]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[30]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8782) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6181 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6364) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6069) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5881);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10255 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6433) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6532) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6260);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049 = ((!N30250) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9684) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9880) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9973) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8814} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8696} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9758};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10183);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9107} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8784} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9451};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481 = !((N30297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437) | ((!N30297) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9481) & N30306));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10065) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9782) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10232} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9605};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10182} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9207} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9977};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10202, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9846} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9296} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9729} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10054};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830} = {1'B0, N26766} + {1'B0, N26768} + {1'B0, N29464};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8758, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10092} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9789} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9565} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10295};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9752) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550 = !((N30297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055) | ((!N30297) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9550) & N30306));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9437);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614 = !((N30297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716) | ((!N30297) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9614) & N30306));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8956} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8985} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9488};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9873} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10012} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10042};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9370} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9824} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8841} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9027};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9848) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9825);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9755} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9213} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10154};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9361);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10239) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10155) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[42]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10033) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9651) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10125) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9068} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9368} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10294};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9905} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9247} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10008};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9497, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9105} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8991} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9761} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9335};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861} = {1'B0, N26750} + {1'B0, N26752} + {1'B0, N29460};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585} = {1'B0, N29466} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9231} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8830};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9195} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9551} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9962};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7984;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7860;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7526) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7654);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7872;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7836)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7960);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8089) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7679;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7776 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7997;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[20] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7995;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9153 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9092 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[21];
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10252} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8942} + {1'B0, N30224};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9049} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9245} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9672};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8649} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10179} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8689};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9380) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8990) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7562 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7923) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[22] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8012 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7602;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193 = !(N29392 | N28088);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9193 | N27939;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9211) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8797} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8966};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9537} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9400} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9597};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8661} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10144} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9169};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[29], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[28]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9563} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10293} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9360};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6620 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5977) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6158) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6346);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[11] = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5859 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6510));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491} = {1'B0, N23050} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[29]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[29]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9516) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9278) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10305} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10006};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8898) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9112) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966 = (!N27939) | (N29392 & N28088);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9966;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 = (!N29392) ^ N28088;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8707) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9769} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9581} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9393};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6279 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6629) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5989) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6168);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9517 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5867) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6519) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6351);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6660 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6324 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6491) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5837) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6211);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9894 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6565) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6026) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6385);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270 = ((!N30248) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9401);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10094) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10184) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8759));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9813) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8989} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9941} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9644};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9717) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9908) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10000) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8848} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8727} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9793};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9408} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9062} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9831} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8876};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8789, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10124} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9598} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9794} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8663};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881} = {1'B0, N26704} + {1'B0, N29452} + {1'B0, N29458};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623} = {1'B0, N29462} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8861} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10237};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7944);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[18] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7909 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7753;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001 = !(N28313 & (!N28113));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9994} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9585} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9270} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10282} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8978};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031 = ((!N30242) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30250));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10031} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9711} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9280};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8837) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9053) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8654) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10131} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9959} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9778};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8721} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9441} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9024};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9974} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10153} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9175};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9446) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9145} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9407} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9205};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[28], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[27]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9367} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10120} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9940};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6472;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6255 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6111) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6393) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6297);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[10] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6005 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6367) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5929));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212} = {1'B0, N23008} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[28]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[28]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9346) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9953} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10128} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10040};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8755) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9192} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9011} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9321};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9178) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017 = (!N28088) | (N28287 & N30226);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9017;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 = (!N28287) ^ N30226;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10228) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9412) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8833} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9383} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9572};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8745} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9480} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9059};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10188} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9792} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9215};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[27], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[26]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8988} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9950} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9760};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6063) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6526) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5876) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6253);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[9] = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5960 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6426));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942} = {1'B0, N22949} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[27]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[27]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6230) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6586) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5940);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9125 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6661) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6121) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6309);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241 = ((!N30246) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10285) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10241} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8650} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10172};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9648) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9246) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10061) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682 = !((N30297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038) | ((!N30297) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9682) & N30306));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9780) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9099} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9404} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10048};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8716);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8812} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9203};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9055);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9876) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9969} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9683} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9252};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9866} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8884} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9674};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8816, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10156} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9638} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8692} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8850};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143} = {1'B0, N26228} + {1'B0, N26230} + {1'B0, N29450};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9219 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7572 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8070;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899} = {1'B0, N30232} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9533} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9881};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6375 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6047) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6503) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6105);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6646) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6465) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6071);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6535 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8774 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5884 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19025);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498 = ((!N30240) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30246));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9623} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9268} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9498};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9477) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9013} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9003} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9183};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9762} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9748} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8778};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8809) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9021) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9715) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8827} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8676} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9375};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9520} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10075} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9093};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10223} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9829} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9251};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[26], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[25]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8815} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9980} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9567};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5948 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6319) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6673) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6488;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[8] = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6558 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6023) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6203;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294} = {1'B0, N23035} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[26]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[26]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8677) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381 = !N30226;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 = !N28313;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133 = !(N30268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10133) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9939) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749 = !((N30297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670) | ((!N30297) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9749) & N30306));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9292} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8882} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8750};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10189} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8660} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8728};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9607, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8723} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9444} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9647};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179} = {1'B0, N26252} + {1'B0, N26254} + {1'B0, N26256};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034 = !(N30232 | N23556);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10034} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9571} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9143};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6419 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6056) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6601) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10108 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5955 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6030) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6139) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6328);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761 = ((!N30234) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30240));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10271} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8899} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8761};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9628} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9815} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10029};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9080) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9314) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8865) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8670} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10164} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9992};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9781} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9356} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8803};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9548) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9777) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8820} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8680} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8996};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9558} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10111} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9129};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10257} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9864} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9288};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[25], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[24]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8847} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10013} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9604};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5932);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5895 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6271) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6622) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6444;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6245) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[7] = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6514 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5982) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6161;
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022} = {1'B0, N22939} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[25]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[25]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9142) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9378) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8926) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9984} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9805} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9619};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8730) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30266) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30268));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10196) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272 = !(N30232 | N23859);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10123) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10030) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9845) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9828} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9025} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9681};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9454} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9482} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10226};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8668, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9982} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8697} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10190} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9217};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951} = {1'B0, N29622} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9272} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9179};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6650) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6054) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6019) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6666) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6377);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6314;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6553) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6432);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9745 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6282) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6196) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5903);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731 = ((!N30238) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30234));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10301} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9917} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9731};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9236} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9427} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9305};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9047} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9818} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9395};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9610) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9841) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10158} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9663} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8665};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8838} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10139} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9164};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10287} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9899} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9328};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[24], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[23]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8883} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10047} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9643};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6578;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5933;
assign N30368 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112 = !N30368;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6112;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5875);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5848 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6223) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6037) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6397);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[6] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6474 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6655) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6010) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6302);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381} = {1'B0, N22929} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[24]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[24]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9206) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9443) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8987) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9609} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9419} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9228};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8781) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30264) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30266));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10259) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245 = !(N30232 | N23861);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9906) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10038);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10093) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10175} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9287} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9442};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9435);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9945) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10217) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10298));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10181) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9998) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810 = !((N30296 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277) | ((!N30296) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9810) & N30305));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10224} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8690} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10080};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9840} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9975} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9263} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10023};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9417, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9035} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10197} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9254} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10015};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000} = {1'B0, N29472} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10245} + {1'B0, N29620};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6262) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6590) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6138 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5971) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5976 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6344) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6508) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5857);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9352 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6045 | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957 = ((!N30236) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30238));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9379} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9951} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8957};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8868} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9045} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9341};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10062} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9081} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8711};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9679) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9902) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9798} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8930} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9979};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9856} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9431} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10174};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9593} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9933} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8657};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[23], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[22]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8916} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10082} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9680};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6643 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5879;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6376 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5998) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6530) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6362);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[5] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6429 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5966) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6067));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094} = {1'B0, N23018} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[23]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[23]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9513) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9220} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9036} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8860};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8834) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30262) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30264));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8651) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501 = !(N30232 | N24239);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10147) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10057) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874 = !((N30296 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907) | ((!N30296) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9874) & N30305));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9865} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9060} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9719};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9968) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8687} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9430} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8917};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8863} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9625} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8892};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9227, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8857} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10049} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9069} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9042};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802} = {1'B0, N26646} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9501} + {1'B0, N29470};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6507) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6147);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6039 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5926) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6606 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6572) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6110) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6471);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8975 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6186) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6296) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947 = ((!N30230) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30236));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10163} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9000} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9947};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10207} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8709} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10130};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10100} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9113} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9697};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9747) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9965) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9411} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8963} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9603};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9887} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8740} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9465};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8870} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9202} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9631};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[22], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[21]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8947} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9362} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9718};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6072 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6600) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5909);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6052) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5866);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6571) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5956 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6064) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5961) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6415);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[4] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6209 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6323) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6596));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458} = {1'B0, N22989} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[22]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[22]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9806) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30258) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30260));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8751) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5993;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5873 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6268 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6674);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6430) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6120) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6244);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5856) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6336) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6173 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6358) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6524) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6424;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6545);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10310 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6061 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5958) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6252);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173 = ((!N30228) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9343)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965) & (!N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935 = !((N30296 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248) | ((!N30296) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9935) & N30305));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9277);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10119) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8712} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9329} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9479};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9470);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9790) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10246) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10148));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10007} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9972} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10203};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9811, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9426} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9657} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8681} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8705};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615} = {1'B0, N27100} + {1'B0, N27102} + {1'B0, N29448};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734 = !(N25457 | N24248);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10212) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10028) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8907);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995 = !((N30296 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888) | ((!N30296) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9995) & N30305));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10213} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9664} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8946};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10258} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8720} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9337};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9397, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9015} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9234} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8986} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9996};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169} = {1'B0, N29398} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9734} + {1'B0, N29446};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763 = !(N30232 | N24241);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8763} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8832} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9615};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9988} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9802} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9008};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9173} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9464} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8826};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9029} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9767} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9958};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30260) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30262));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8704) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8894) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9188} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9851} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10025};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9151} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8938} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9735};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9342) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9577) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9109) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8853} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8700} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10200};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9924} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8765} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9505};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8905} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10211} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9669};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[21], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[20]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9970} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8685} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8984};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6416 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6070);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6015;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6191;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5897 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6180);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6371;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6080);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6192);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5863 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6142 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6308) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6118) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6480);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[3] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6085 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6278) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6450) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5899);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178} = {1'B0, N22959} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[21]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[21]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9174) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9409) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8965 | N30228);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30256) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30258));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8805) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8675} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10149} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9076};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10016} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9842} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9776};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9742} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10279} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9543};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10024) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9645) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8953) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9871) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9661} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10193} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8695};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9210} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8795} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8974};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9705} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8743} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10247};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[20], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[19]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9241} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8715} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10001};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6370 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6050) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5850);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6029 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6613;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6551 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6470);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5954 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6014) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6455);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6665 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6208) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6626);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5883 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6434) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6263) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6150);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[2] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6341 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5852) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5972));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906} = {1'B0, N22969} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[20]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[20]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10086) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9712) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9018) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9932) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9267} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9833} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10010};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8843} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9579} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8800};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9244) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9474) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10178) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10090) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9512);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9632) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10003));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9897} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9094} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10041};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9757, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9364} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10095} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9594} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8658};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960 = !(N30232 | N24250);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784} = {1'B0, N26726} + {1'B0, N29396} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8960};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30254) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30256));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8862) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10143} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10169} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8736};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9649} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9458} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9589};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9552} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10308} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9351};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8773} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9315} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9514};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[19], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9276} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9473} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10037};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6476) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6411) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5919;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5916) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6388) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6124) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6213);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6164 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6136) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6225);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6104;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6151) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5914);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6383 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6518) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6386);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6202) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6425 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6327) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5839) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6494);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[1] = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6645 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6567) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6001) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6464);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259} = {1'B0, N22979} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[19]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[19]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6490) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6533) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6027);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5889) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5920) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6583);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5992;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6162 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6126) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6461);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6326 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5981) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5938) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6404);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6563 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5925) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6096) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6580);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6598 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6321) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6291) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6338);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6090 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6454) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6631) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6170);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[0] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6520 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6055) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N6354));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10142) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9772) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9077) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9993) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8893} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9448} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9640};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10187} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9389} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8652};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9310) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9544) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10145) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10248);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10242) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8897} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9521} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8746};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9108, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8760} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10215} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8958} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9730};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949 = !(N30232 | N24268);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117} = {1'B0, N26742} + {1'B0, N26744} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9949};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30244) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30254));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8923) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8785} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9784} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10060};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9258} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9071} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9167};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9359} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10135} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9160};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10284} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10106} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9324};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[18], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10070} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10253} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9087};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989} = {1'B0, N23378} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[18]};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10205) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9837) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9140) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10053) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10236} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9066} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9249};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9827} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9198} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9936};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9439) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9676) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116 = !((N30296 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115) | ((!N30296) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10116) & N30305));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10064} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9882} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9934};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055 = !((N30295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507) | ((!N30295) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9888));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10055) & N30304));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9243, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8872} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10288} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9374} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9858};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177 = !(N30232 | N24653);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499} = {1'B0, N26734} + {1'B0, N26736} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9177};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9549);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9467) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10299) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9857));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10209) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176 = !((N30295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766) | ((!N30295) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10176) & N30304));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10269) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9106} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9557} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8777};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10127, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9130} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10074} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10039};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152 = !(N30232 | N24633);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633} = {1'B0, N27092} + {1'B0, N27094} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10152};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30250) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30252));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9046) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10005} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9499} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9300};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10227} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10052} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8901};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9898) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30250));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9204) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10115) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9879} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8725} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8879};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10265} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9298} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9562};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8980} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9750} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8752};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9608) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9372) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8817} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8886} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8729};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8908);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9952) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10266) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10302));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30252) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30244));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8983) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9884} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10117} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9694};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9529} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9438} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8806};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8950} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9964} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9722};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10114} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9930} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9131};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8943} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9901} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9714};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9123} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10076} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9893};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12310);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9115);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238 = !((N30295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101) | ((!N30295) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10238) & N30304));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9918} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10091} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9165};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9586);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9306) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8662) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9698));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297 = !((N30295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736) | ((!N30295) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10297) & N30304));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8766);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10101);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736 | N30295);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9144) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8686) & N30304));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9476} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[2]} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10296} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10138};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9030} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9336} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8804} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9863};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9344} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10112} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10304} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9410};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8717} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8968} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9671} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9737};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9147, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8791} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8995} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9764} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9057};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30242) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N24635));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9104) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688} = {1'B0, N29618} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9633} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8928};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10020) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30248));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9339) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9804) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9103} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9678} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9485};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9022} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10240} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9791};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9910} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8924} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9432};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9961) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8693} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9494} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10046};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9707);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9795) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10173) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10157));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9744) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9508) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9870} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10220} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9686};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9136} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9665} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8713};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10290} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10056} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9330};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9074} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10085} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9101};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9492} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8780} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9524};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405 = !(N30232 | N30250);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30248) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30242));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9170) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9405} + {1'B0, N29616} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10268};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9573) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9293} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9920} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8688};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8813} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9269} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10032};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9691} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10177} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8735};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9641) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9868) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691 = !(N30232 | N24662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30246) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N24642));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9240) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440} = {1'B0, N27231} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8691} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9912};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9097} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8921} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9826};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30240) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30246));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9406) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8775);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9639) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10081) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10009));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10219} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8757} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9285};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8932} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9701} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9403};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9048} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9566} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9820};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9931) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9471) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9708) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10088} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8749} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10262};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9536} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8845} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10274};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10150} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8741} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9172};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635 = !(N30232 | N24642);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N25288) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N24644));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9304) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104} = {1'B0, N27456} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9635} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9532};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30234));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9542) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9555);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9475) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9989) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9861));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10071} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9725} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10078};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8767} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9440} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9510};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9308} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9602} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10066};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874 = !(N30232 | N30246);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30234) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30240));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9369) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797} = {1'B0, N27448} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8874} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9139};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9770) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9903} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10160} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10104};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10250} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10186} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9209};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9834) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30236) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30238));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9606) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859 = !(N30232 | N30240);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N30238) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N25313));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9436) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222} = {1'B0, N27640} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9859} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8786};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9334} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9527} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8878};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9182} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9117} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9889};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30230) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9673) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8655);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9317) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9895) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9706));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9925} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8952} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9133};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9797} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9642} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8819};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084 = !(N30232 | N30234);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9564 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N7975 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9736);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N25297) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N25295));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9504) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710} = {1'B0, N27844} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9084} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10122};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069 = !(N30232 | N30238);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N25852) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N30236));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9570) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10069} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9759};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402 & N30228) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402) & N30230));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741 & N30224) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9741) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10292} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10281} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9710};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10072} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10222} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9090};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9402);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801 & N29556) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9801) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311 = !(N30232 | N30236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669 & N25854) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669) & N25852));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9637) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9311} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9366};
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9768} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9942} + {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9546};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277 = !(N30232 | N30230);
assign {DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2], DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[1]} = {1'B0, DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N10277} + {1'B0, N30226};
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704 = !(N30228 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N8669);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[1] = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9001) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9704) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N9381));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[1] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12230) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12278)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[2]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[2]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[3] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12112 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12509) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12376);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12151) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11958)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[4]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[4]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12346 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12432) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12291);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12069) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12101)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[6]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[6]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[7] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12421 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12350) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12207);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11996) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12083)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[8]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[8]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[9] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12320 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12270) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12128);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11915) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11920)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[10]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[10]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[11] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12061 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12185) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12052);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12467) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12210)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[12]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[12]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[13] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12281 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12104) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11973);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[14] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[15] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12243 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12031) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12519);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12348) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12410)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12266);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[16] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[17] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12161 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11948) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12444);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12220) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12169)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[18]) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11989));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12250 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12148) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12014);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12498) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12192)) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12120) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12259));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12405 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11906);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12044 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12178);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12317 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12458);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11966 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12094);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12235 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12381);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12512 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12022);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12155 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12294);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12436 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11942);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12072 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12212);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12354 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12491);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12000 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12132);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12272 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12416);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11919 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12054);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12189 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12329);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12469 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11977);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12108 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12245);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12522 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12164 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12033);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12446 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12305);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182 = !(N29502 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11951);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464 = !(N22618 | N29506);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12008 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12501);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12283 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12140);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12424 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11929);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12059 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12197);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12415 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12298 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12355) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12255);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12337 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12476);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11984 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12117);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12246 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12400 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12330 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302 = (N29510 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12391) | N21795;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12302;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12443 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12356);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107 = N29679 & N29681;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156 = N22305 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273 = N21999 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11983;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12057;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12137;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12007 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12423) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12279;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11925 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12333) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12196;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12473 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464 & N22305) | N22309;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024 & N21999) | N22003;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11976 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11921) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12418;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12107) | N20660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12160) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12030;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12217) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12076;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[48] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12133) ^ N20538;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & N20492) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[48];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219 | N18660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470 = N29667 & N29669;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999 = N21993 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12515;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12045;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12202;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12371;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12524;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11981) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12472;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12397 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12449) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12308;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12226 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12286) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12146;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12063 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12123) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11991;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11910 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11968) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12460;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12383 & N21993) | N21988;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12328 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12214 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12276) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12135;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12470) | N21782;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12518) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12387;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11945) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12440;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11901 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12005 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12497));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[47] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12494 ^ N21075;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[47];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12188 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12075;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12236;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242 = N21765 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12406;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11933;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12084;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12249;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12331) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12194;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12110 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12168) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12036;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11956 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12013) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12504;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12427 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12481) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12344;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12261 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12321) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12180;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12099 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12156) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12024;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12055 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11944 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12002) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12495;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211 & N21765) | N21769;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12242) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12103;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12299) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12157;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12115 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12357 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12218));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[46] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12213 ^ N21090;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[46];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972 = N29566 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12073;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12404;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12082;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11953 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11931) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12426;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12258 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12234) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12095;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11941 & N29566) | N29510;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11972) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12466;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12027) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12516;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12335 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12077 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11946));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[45] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11943 ^ N21080;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[45];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12435;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12121;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12448;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12307 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12285) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12143;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11988 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11965) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12457;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12295 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12273) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12131;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12324) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12184;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12384) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12239;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11927 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12441 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12300));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[44] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12297 ^ N21085;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[44];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12154;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12479;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12011) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12503;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12341 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12318) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12177;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12021 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11999) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12492;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12051) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11914;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12100) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11969;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12138 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12158 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12028));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[43] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12023 ^ N21070;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[43];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12513;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12201;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12367) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12225;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12062 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12043) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11907;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12380 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12353) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12211;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12411) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12269;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12463) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12322;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12362 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12517 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12385));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[42] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12382 ^ N21100;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[42];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12453;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12313 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12127) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11995;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12181) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12047;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11950 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12240 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12102));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[41] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12097 ^ N21105;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[41];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12174;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12040 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12487) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12349;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12364 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11911) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12407;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11970 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12464));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[40] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12459 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12163;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[40];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11902;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12401 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12206) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12068;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12035 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12263) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12125;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12323 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12182));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[39] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12179 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12390;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[39];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12254;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12116 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11937) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12431;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12394 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11992) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12484;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12048 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11912));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[38] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11909 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11975;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[38];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11985;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12475 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12290) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12150;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11923 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12345) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12203;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12408 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12265));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[37] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12260 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12187;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[37];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12336;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12198 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12017) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12508;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12360 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12065) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11935;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12126 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11993));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[36] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11990 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12414;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[36];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12375) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12229);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12485 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12347));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[35] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12264) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11998;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[35];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12090) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11961);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12204 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12066));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[34] = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12124) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12209;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[34];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11936 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12429));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[33] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12373 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12434;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[33];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12288 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12149));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[32] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12086 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12020;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[32];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12015 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12506));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[31] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12450 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12232;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[31];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12374 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12227));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[30] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12171 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12456;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[30];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12087 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11959));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[29] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11898 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12042;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[29];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12451 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12311));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[28] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12251 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12257;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[28];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13351) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13411)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13387);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13354 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13406) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13347);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12172 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12037));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[27] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11928 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12478;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[27];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N11899 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12399));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[26] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12282 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12060;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[26];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13371;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13397 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13355) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13349);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13399 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13380));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13341;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13359 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13407) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13375);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13367 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13392);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13365 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13348));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13391) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13373 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13383);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13339) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13374);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12252 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12113));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[25] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12009 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N12284;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13041 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[25];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13340) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13376);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4] | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13384) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13402);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13393) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13405)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13337);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8] | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13409) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13343);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12] | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13352) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13368);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13362) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13346)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13388);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13379 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13356) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13334);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16] | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13377) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13395);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20] | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13404) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21])) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13398);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13370) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13332)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13358));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541 = ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13360) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386)) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13394);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531 = (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13475) ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13386;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3] = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13470 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N544;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13472 ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N543;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0] = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N541;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0] ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N542;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[22]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13492 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13540 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13490 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13591 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670 = (N30278 & N18886) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N701);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185 = !(a_exp[7] & a_exp[0]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047 = !((a_exp[6] & a_exp[5]) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13187);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13185 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19047);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N19054;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225 = !(((a_man[0] | a_man[1]) | a_man[2]) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13221);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208 = !(a_man[10] | a_man[9]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227 = !(a_man[6] | a_man[5]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216 = !(a_man[8] | a_man[7]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236 = !(N30313 | a_man[3]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13208 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13227) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13216) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13236);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13225) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13219) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13230) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13240);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__19 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__24;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288 = ((a_exp[7] | a_exp[6]) | a_exp[0]) | a_exp[5];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292 = ((a_exp[4] | a_exp[2]) | a_exp[3]) | a_exp[1];
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13288 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13292);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487 = DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__17 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__68) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[22] = (N30273 & N30270) | ((!N30273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N670);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[11]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[10]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[13]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[12]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[7]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[6]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[9]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[8]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[19]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[18]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[21]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[20]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13612 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[15]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[14]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[17]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[16]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13511 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13610 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[3]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[2]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[5]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[4]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555 = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[1]) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[0]);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13558 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669 = (N30281 & N18971) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N700);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[21] = (N30272 & N30270) | ((!N30272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13548 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13617 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13571 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13635 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13512 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13577 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13527 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13598 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13628 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13576 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13589 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13503 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13639 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13522 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668 = (N30279 & N19020) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N699);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[20] = (N30273 & N30270) | ((!N30273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13518 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13583 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13534 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13604 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13629 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13541 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13497 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13565 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13596 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13539 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13555 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13609) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13623 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13491 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667 = (N30282 & N19000) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N698);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[19] = (N30276 & N30270) | ((!N30276) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13603 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13621 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13563 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13582 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13510 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13638);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13611 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666 = (N30282 & N19030) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N697);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[18] = (N30274 & N30270) | ((!N30274) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13570 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13587 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13526 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13547 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13627 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13574);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13578 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665 = (N30279 & N19010) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N696);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[17] = (N30275 & N30270) | ((!N30275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13533 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13554 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13496 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13517 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13595 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13507);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13542 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664 = (N30281 & N18990) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N695);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[16] = (N30274 & N30270) | ((!N30274) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13502 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13521 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13616 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13634 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13566));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13562 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13513);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663 = (N30283 & N19040) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N694);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[15] = (N30275 & N30270) | ((!N30275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13569 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13525 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13630);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662 = (N30278 & N19050) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N693);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[14] = (N30274 & N30270) | ((!N30274) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13532 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13495 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13597);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661 = (N30280 & N19099) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N692);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[13] = (N30275 & N30270) | ((!N30275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13501 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13615 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13564);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660 = (N30278 & N19109) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N691);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[12] = (N30272 & N30270) | ((!N30272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13553 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13581 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13528);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659 = (N30284 & N19119) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N690);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[11] = (N30272 & N30270) | ((!N30272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13608 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13546 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13498);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658 = (N30278 & N19149) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N689);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[10] = (N30275 & N30270) | ((!N30275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13506 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13516 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13618);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657 = (N30280 & N19060) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N688);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[9] = (N30274 & N30270) | ((!N30274) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13560 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[3]) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13633 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13584);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656 = (N30283 & N19129) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N687);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[8] = (N30272 & N30270) | ((!N30272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13602 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13588);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655 = (N30280 & N19159) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N686);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[7] = (N30273 & N30270) | ((!N30273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13605);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654 = (N30283 & N19139) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N685);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[6] = (N30276 & N30270) | ((!N30276) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13535);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653 = (N30282 & N19070) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N684);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[5] = (N30273 & N30270) | ((!N30273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13622);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652 = (N30281 & N19080) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N683);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[4] = (N30273 & N30270) | ((!N30273) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13556);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651 = (N30282 & N19233) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N682);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[3] = (N30276 & N30270) | ((!N30276) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650 = (N30281 & N19223) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N681);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[2] = (N30275 & N30270) | ((!N30275) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13575);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649 = (N30280 & N19275) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N680);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[1] = (N30274 & N30270) | ((!N30274) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13545 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13509);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648 = (N30279 & N19410) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N679);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[0] = (N30272 & N30270) | ((!N30272) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647 = a_exp[7] & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N639;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N487 & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__82));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N759;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026 = !DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14019;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[30] = (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N580) | ((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N14026) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N647);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__219 & (!N30278));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863 = !((N30281 & N20175) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13863);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[29] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818 = !((N30280 & N20182) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13818);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[28] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877 = !((N30283 & N19891) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13531));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13877);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[27] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832 = !((N30283 & N19768) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13551));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13832);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[26] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786 = !((N30279 & N19900) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13549));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13786);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[25] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845 = !((N30279 & N19909) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13594));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13845);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[24] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800 = !((N30282 & N20144) | (DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13822 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13601));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13809 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13800);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[23] = (N18835 & N18839) | ((!N18835) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5515 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5409);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[5] | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N5424);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N577 = a_sign ^ DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N757;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N667 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N665) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N668) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N666;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N653 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N652) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N663);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N651 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N655) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N658);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947 = ((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N659 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N656) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N661) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N660;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13937) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N669) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13947) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N664);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925 = ((N19633 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N645) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N646) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N640;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13925 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N641) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N642);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969 = !(DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N643 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N644);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939 = !((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13969 & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13957) & (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N648));
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955 = !(((DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N649 | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N650) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13939) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N654);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934 = !(((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13955) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N657) | DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N662);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578 = !((((!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13970) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13943) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13940) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N13934);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579 = !((((!N18881) | (!DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N578)) | N18678) | N18879);
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[31] = (N30284 & N18664) | ((!N30284) & DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_N579);
reg x_reg_L0_30__I3803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_30__I3803_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[30];
	end
assign N9100 = x_reg_L0_30__I3803_QOUT;
reg x_reg_L1_0__I3805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__I3805_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[0];
	end
assign x[0] = x_reg_L1_0__I3805_QOUT;
reg x_reg_L1_1__I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__I3806_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[1];
	end
assign x[1] = x_reg_L1_1__I3806_QOUT;
reg x_reg_L1_2__I3807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__I3807_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[2];
	end
assign x[2] = x_reg_L1_2__I3807_QOUT;
reg x_reg_L1_3__I3808_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__I3808_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[3];
	end
assign x[3] = x_reg_L1_3__I3808_QOUT;
reg x_reg_L1_4__I3809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__I3809_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[4];
	end
assign x[4] = x_reg_L1_4__I3809_QOUT;
reg x_reg_L1_5__I3810_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__I3810_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[5];
	end
assign x[5] = x_reg_L1_5__I3810_QOUT;
reg x_reg_L1_6__I3811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__I3811_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[6];
	end
assign x[6] = x_reg_L1_6__I3811_QOUT;
reg x_reg_L1_7__I3812_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__I3812_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[7];
	end
assign x[7] = x_reg_L1_7__I3812_QOUT;
reg x_reg_L1_8__I3813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__I3813_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[8];
	end
assign x[8] = x_reg_L1_8__I3813_QOUT;
reg x_reg_L1_9__I3814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__I3814_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[9];
	end
assign x[9] = x_reg_L1_9__I3814_QOUT;
reg x_reg_L1_10__I3815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__I3815_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[10];
	end
assign x[10] = x_reg_L1_10__I3815_QOUT;
reg x_reg_L1_11__I3816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__I3816_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[11];
	end
assign x[11] = x_reg_L1_11__I3816_QOUT;
reg x_reg_L1_12__I3817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__I3817_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[12];
	end
assign x[12] = x_reg_L1_12__I3817_QOUT;
reg x_reg_L1_13__I3818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__I3818_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[13];
	end
assign x[13] = x_reg_L1_13__I3818_QOUT;
reg x_reg_L1_14__I3819_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__I3819_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[14];
	end
assign x[14] = x_reg_L1_14__I3819_QOUT;
reg x_reg_L1_15__I3820_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__I3820_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[15];
	end
assign x[15] = x_reg_L1_15__I3820_QOUT;
reg x_reg_L1_16__I3821_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__I3821_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[16];
	end
assign x[16] = x_reg_L1_16__I3821_QOUT;
reg x_reg_L1_17__I3822_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__I3822_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[17];
	end
assign x[17] = x_reg_L1_17__I3822_QOUT;
reg x_reg_L1_18__I3823_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__I3823_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[18];
	end
assign x[18] = x_reg_L1_18__I3823_QOUT;
reg x_reg_L1_19__I3824_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__I3824_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[19];
	end
assign x[19] = x_reg_L1_19__I3824_QOUT;
reg x_reg_L1_20__I3825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__I3825_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[20];
	end
assign x[20] = x_reg_L1_20__I3825_QOUT;
reg x_reg_L1_21__I3826_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__I3826_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[21];
	end
assign x[21] = x_reg_L1_21__I3826_QOUT;
reg x_reg_L1_22__I3827_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__I3827_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[22];
	end
assign x[22] = x_reg_L1_22__I3827_QOUT;
reg x_reg_L1_23__I3828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__I3828_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[23];
	end
assign x[23] = x_reg_L1_23__I3828_QOUT;
reg x_reg_L1_24__I3829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__I3829_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[24];
	end
assign x[24] = x_reg_L1_24__I3829_QOUT;
reg x_reg_L1_25__I3830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__I3830_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[25];
	end
assign x[25] = x_reg_L1_25__I3830_QOUT;
reg x_reg_L1_26__I3831_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__I3831_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[26];
	end
assign x[26] = x_reg_L1_26__I3831_QOUT;
reg x_reg_L1_27__I3832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__I3832_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[27];
	end
assign x[27] = x_reg_L1_27__I3832_QOUT;
reg x_reg_L1_28__I3833_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__I3833_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[28];
	end
assign x[28] = x_reg_L1_28__I3833_QOUT;
reg x_reg_L1_29__I3834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__I3834_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[29];
	end
assign x[29] = x_reg_L1_29__I3834_QOUT;
reg x_reg_L1_30__I3835_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__I3835_QOUT <= N9100;
	end
assign x[30] = x_reg_L1_30__I3835_QOUT;
reg x_reg_L1_31__I3836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I3836_QOUT <= DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I3836_QOUT;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[32] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[33] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[34] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[35] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_x[36] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__42[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__61[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__195[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__198[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[3] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[4] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[5] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[6] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[7] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[8] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[9] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[10] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[11] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[12] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[13] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[14] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[15] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[16] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[17] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[18] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[19] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[20] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[21] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[22] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__201[49] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W0[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[0] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[43] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[44] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[45] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__203__W1[46] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[23] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[24] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[25] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[26] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[27] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[28] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[29] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__210[30] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[1] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[2] = 1'B0;
assign DFT_compute_cynw_cm_float_sin_E8_M23_2_inst_inst_cellmath__215[4] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  urP1TQHarh9B : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



