/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:20:26 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_sin_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__66,
	inst_cellmath__67,
	inst_cellmath__68,
	inst_cellmath__69,
	inst_cellmath__82;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__200,
	inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire  inst_cellmath__219;
wire N487,N541,N542,N543,N544,N545,N577 
	,N578,N579,N580,N582,N583,N584,N585,N586 
	,N587,N588,N589,N590,N591,N592,N593,N594 
	,N595,N596,N597,N598,N599,N600,N601,N602 
	,N603,N604,N605,N606,N607,N608,N609,N610 
	,N611,N612,N613,N614,N615,N616,N617,N618 
	,N619,N620,N621,N622,N623,N624,N625,N626 
	,N627,N628,N629,N630,N631,N632,N633,N634 
	,N635,N636,N637,N639,N640,N641,N642,N643 
	,N644,N645,N646,N647,N648,N649,N650,N651 
	,N652,N653,N654,N655,N656,N657,N658,N659 
	,N660,N661,N662,N663,N664,N665,N666,N667 
	,N668,N670,N671,N672,N673,N674,N675,N676 
	,N677,N679,N680,N681,N682,N683,N684,N685 
	,N686,N687,N688,N689,N690,N691,N692,N693 
	,N694,N695,N696,N697,N698,N699,N700,N701 
	,N733,N734,N735,N736,N737,N738,N739,N740 
	,N741,N742,N743,N744,N745,N746,N747,N748 
	,N749,N750,N751,N752,N753,N754,N755,N756 
	,N757,N759,N760,N761,N762,N763,N764,N765 
	,N766,N767,N768,N769,N770,N771,N772,N773 
	,N774,N775,N776,N777,N778,N779,N780,N781 
	,N782,N3584,N3657,N3658,N3659,N3660,N3661,N3662 
	,N3665,N3666;
cynw_cm_float_sin_inst_blk01_cellmath__39_bdw1946085813_bdw cynw_cm_float_sin_I0 (.inst_blk01_cellmath__39_out0({N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582}), .inst_blk01_cellmath__39_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_sin_inst_cellmath__42_0_bdw1946085813_bdw cynw_cm_float_sin_I1 (.inst_cellmath__42_0_out0({inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__42_0_in0({a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_sin_inst_cellmath__48_bdw1946085813_bdw cynw_cm_float_sin_I2 (.inst_cellmath__48_out0({N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733}), .inst_cellmath__48_in0({inst_cellmath__42[5], inst_cellmath__42[4], inst_cellmath__42[3], inst_cellmath__42[2], inst_cellmath__42[1], inst_cellmath__42[0]}), .inst_cellmath__48_in1({N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608}));
cynw_cm_float_sin_inst_cellmath__61_0_bdw1946085813_bdw cynw_cm_float_sin_I3 (.inst_cellmath__61_0_out0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17], inst_cellmath__61[16], inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__61_0_in0({N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733}));
INVXL cynw_cm_float_sin_I296 (.Y(N3657), .A(inst_cellmath__61[10]));
INVXL cynw_cm_float_sin_I297 (.Y(N3658), .A(N3657));
INVXL cynw_cm_float_sin_I298 (.Y(N3659), .A(inst_cellmath__61[6]));
INVXL cynw_cm_float_sin_I299 (.Y(N3660), .A(N3659));
INVXL cynw_cm_float_sin_I300 (.Y(N3661), .A(inst_cellmath__61[2]));
INVXL cynw_cm_float_sin_I301 (.Y(N3662), .A(N3661));
INVXL cynw_cm_float_sin_I304 (.Y(N3665), .A(inst_cellmath__61[8]));
INVXL cynw_cm_float_sin_I305 (.Y(N3666), .A(N3665));
INVXL cynw_cm_float_sin_I4 (.Y(inst_cellmath__115__W1[0]), .A(inst_cellmath__61[16]));
cynw_cm_float_sin_inst_cellmath__195__80__2WWMM_2WWMM_bdw1946085813_bdw cynw_cm_float_sin_I5 (.inst_cellmath__195__80__2WWMM_2WWMM_out0({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0], inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0], N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760}), .inst_cellmath__195__80__2WWMM_2WWMM_in0({inst_cellmath__61[22], inst_cellmath__61[21], inst_cellmath__61[20], inst_cellmath__61[19], inst_cellmath__61[18], inst_cellmath__61[17]}));
cynw_cm_float_sin_inst_cellmath__198_0_bdw1946085813_bdw cynw_cm_float_sin_I6 (.inst_cellmath__198_0_out0({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17], inst_cellmath__198[16], inst_cellmath__198[15], inst_cellmath__198[14], inst_cellmath__198[13], inst_cellmath__198[12], inst_cellmath__198[11], inst_cellmath__198[10], inst_cellmath__198[9], inst_cellmath__198[8], inst_cellmath__198[7], inst_cellmath__198[6], inst_cellmath__198[5], inst_cellmath__198[4], inst_cellmath__198[3], inst_cellmath__198[2], inst_cellmath__198[1], inst_cellmath__198[0]}), .inst_cellmath__198_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], inst_cellmath__61[10], inst_cellmath__61[9], inst_cellmath__61[8], inst_cellmath__61[7], inst_cellmath__61[6], inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], inst_cellmath__61[2], inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__198_0_in1({inst_cellmath__115__W1[0]}));
cynw_cm_float_sin_inst_cellmath__203_0_bdw1946085813_bdw cynw_cm_float_sin_I7 (.inst_cellmath__203_0_out0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__203_0_out1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__203_0_in0({inst_cellmath__61[15], inst_cellmath__61[14], inst_cellmath__61[13], inst_cellmath__61[12], inst_cellmath__61[11], N3658, inst_cellmath__61[9], N3666, inst_cellmath__61[7], N3660, inst_cellmath__61[5], inst_cellmath__61[4], inst_cellmath__61[3], N3662, inst_cellmath__61[1], inst_cellmath__61[0]}), .inst_cellmath__203_0_in1({inst_cellmath__198[32], inst_cellmath__198[31], inst_cellmath__198[30], inst_cellmath__198[29], inst_cellmath__198[28], inst_cellmath__198[27], inst_cellmath__198[26], inst_cellmath__198[25], inst_cellmath__198[24], inst_cellmath__198[23], inst_cellmath__198[22], inst_cellmath__198[21], inst_cellmath__198[20], inst_cellmath__198[19], inst_cellmath__198[18], inst_cellmath__198[17]}), .inst_cellmath__203_0_in2({inst_cellmath__197[19], inst_cellmath__197[18], inst_cellmath__197[17], inst_cellmath__197[16], inst_cellmath__197[15], inst_cellmath__197[14], inst_cellmath__197[13], inst_cellmath__197[12], inst_cellmath__197[11], inst_cellmath__197[10], inst_cellmath__197[9], inst_cellmath__197[8], inst_cellmath__197[7], inst_cellmath__197[6], inst_cellmath__197[5], inst_cellmath__197[4], inst_cellmath__197[3], inst_cellmath__197[2], inst_cellmath__197[1], inst_cellmath__197[0]}), .inst_cellmath__203_0_in3({N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760}), .inst_cellmath__203_0_in4({inst_cellmath__115__W1[0]}));
cynw_cm_float_sin_inst_cellmath__201_0_bdw1946085813_bdw cynw_cm_float_sin_I8 (.inst_cellmath__201_0_out0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}), .inst_cellmath__201_0_in0({inst_cellmath__203__W1[46], inst_cellmath__203__W1[45], inst_cellmath__203__W1[44], inst_cellmath__203__W1[43], inst_cellmath__203__W1[42], inst_cellmath__203__W1[41], inst_cellmath__203__W1[40], inst_cellmath__203__W1[39], inst_cellmath__203__W1[38], inst_cellmath__203__W1[37], inst_cellmath__203__W1[36], inst_cellmath__203__W1[35], inst_cellmath__203__W1[34], inst_cellmath__203__W1[33], inst_cellmath__203__W1[32], inst_cellmath__203__W1[31], inst_cellmath__203__W1[30], inst_cellmath__203__W1[29], inst_cellmath__203__W1[28], inst_cellmath__203__W1[27], inst_cellmath__203__W1[26], inst_cellmath__203__W1[25], inst_cellmath__203__W1[24], inst_cellmath__203__W1[23], inst_cellmath__203__W1[22], inst_cellmath__203__W1[21], inst_cellmath__203__W1[20], inst_cellmath__203__W1[19], inst_cellmath__203__W1[18], inst_cellmath__203__W1[17], inst_cellmath__203__W1[16], inst_cellmath__203__W1[15], inst_cellmath__203__W1[14], inst_cellmath__203__W1[13], inst_cellmath__203__W1[12], inst_cellmath__203__W1[11], inst_cellmath__203__W1[10], inst_cellmath__203__W1[9], inst_cellmath__203__W1[8], inst_cellmath__203__W1[7], inst_cellmath__203__W1[6], inst_cellmath__203__W1[5], inst_cellmath__203__W1[4], inst_cellmath__203__W1[3], inst_cellmath__203__W1[2], inst_cellmath__203__W1[1], inst_cellmath__203__W1[0]}), .inst_cellmath__201_0_in1({inst_cellmath__203__W0[46], inst_cellmath__203__W0[45], inst_cellmath__203__W0[44], inst_cellmath__203__W0[43], inst_cellmath__203__W0[42], inst_cellmath__203__W0[41], inst_cellmath__203__W0[40], inst_cellmath__203__W0[39], inst_cellmath__203__W0[38], inst_cellmath__203__W0[37], inst_cellmath__203__W0[36], inst_cellmath__203__W0[35], inst_cellmath__203__W0[34], inst_cellmath__203__W0[33], inst_cellmath__203__W0[32], inst_cellmath__203__W0[31], inst_cellmath__203__W0[30], inst_cellmath__203__W0[29], inst_cellmath__203__W0[28], inst_cellmath__203__W0[27], inst_cellmath__203__W0[26], inst_cellmath__203__W0[25], inst_cellmath__203__W0[24], inst_cellmath__203__W0[23], inst_cellmath__203__W0[22], inst_cellmath__203__W0[21], inst_cellmath__203__W0[20], inst_cellmath__203__W0[19], inst_cellmath__203__W0[18], inst_cellmath__203__W0[17], inst_cellmath__203__W0[16], inst_cellmath__203__W0[15], inst_cellmath__203__W0[14], inst_cellmath__203__W0[13], inst_cellmath__203__W0[12], inst_cellmath__203__W0[11], inst_cellmath__203__W0[10], inst_cellmath__203__W0[9], inst_cellmath__203__W0[8], inst_cellmath__203__W0[7], inst_cellmath__203__W0[6], inst_cellmath__203__W0[5], inst_cellmath__203__W0[4], inst_cellmath__203__W0[3], inst_cellmath__203__W0[2], inst_cellmath__203__W0[1], inst_cellmath__203__W0[0]}), .inst_cellmath__201_0_in2({inst_cellmath__195[29], inst_cellmath__195[28], inst_cellmath__195[27], inst_cellmath__195[26], inst_cellmath__195[25], inst_cellmath__195[24], inst_cellmath__195[23], inst_cellmath__195[22], inst_cellmath__195[21], inst_cellmath__195[20], inst_cellmath__195[19], inst_cellmath__195[18], inst_cellmath__195[17], inst_cellmath__195[16], inst_cellmath__195[15], inst_cellmath__195[14], inst_cellmath__195[13], inst_cellmath__195[12], inst_cellmath__195[11], inst_cellmath__195[10], inst_cellmath__195[9], inst_cellmath__195[8], inst_cellmath__195[7], inst_cellmath__195[6], inst_cellmath__195[5], inst_cellmath__195[4], inst_cellmath__195[3], inst_cellmath__195[2], inst_cellmath__195[1], inst_cellmath__195[0]}));
cynw_cm_float_sin_inst_cellmath__200_0_bdw1946085813_bdw cynw_cm_float_sin_I9 (.inst_cellmath__200_0_out0({inst_cellmath__200[48], inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0], inst_cellmath__200[24], inst_cellmath__200[23], inst_cellmath__200[22], inst_cellmath__200[21], inst_cellmath__200[20], inst_cellmath__200[19], inst_cellmath__200[18], inst_cellmath__200[17], inst_cellmath__200[16], inst_cellmath__200[15], inst_cellmath__200[14], inst_cellmath__200[13], inst_cellmath__200[12], inst_cellmath__200[11], inst_cellmath__200[10], inst_cellmath__200[9], inst_cellmath__200[8], inst_cellmath__200[7], inst_cellmath__200[6], inst_cellmath__200[5], inst_cellmath__200[4], inst_cellmath__200[3], inst_cellmath__200[2], inst_cellmath__200[1], inst_cellmath__200[0]}), .inst_cellmath__200_0_in0({inst_cellmath__201[49], inst_cellmath__201[48], inst_cellmath__201[47], inst_cellmath__201[46], inst_cellmath__201[45], inst_cellmath__201[44], inst_cellmath__201[43], inst_cellmath__201[42], inst_cellmath__201[41], inst_cellmath__201[40], inst_cellmath__201[39], inst_cellmath__201[38], inst_cellmath__201[37], inst_cellmath__201[36], inst_cellmath__201[35], inst_cellmath__201[34], inst_cellmath__201[33], inst_cellmath__201[32], inst_cellmath__201[31], inst_cellmath__201[30], inst_cellmath__201[29], inst_cellmath__201[28], inst_cellmath__201[27], inst_cellmath__201[26], inst_cellmath__201[25], inst_cellmath__201[24], inst_cellmath__201[23], inst_cellmath__201[22], inst_cellmath__201[21], inst_cellmath__201[20], inst_cellmath__201[19], inst_cellmath__201[18], inst_cellmath__201[17], inst_cellmath__201[16], inst_cellmath__201[15], inst_cellmath__201[14], inst_cellmath__201[13], inst_cellmath__201[12], inst_cellmath__201[11], inst_cellmath__201[10], inst_cellmath__201[9], inst_cellmath__201[8], inst_cellmath__201[7], inst_cellmath__201[6], inst_cellmath__201[5], inst_cellmath__201[4], inst_cellmath__201[3], inst_cellmath__201[2], inst_cellmath__201[1], inst_cellmath__201[0]}));
cynw_cm_float_sin_inst_cellmath__19_0_bdw1946085813_bdw cynw_cm_float_sin_I10 (.inst_cellmath__19_0_out0(inst_cellmath__19), .inst_cellmath__19_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_sin_inst_cellmath__24_0_bdw1946085813_bdw cynw_cm_float_sin_I11 (.inst_cellmath__24_0_out0(inst_cellmath__24), .inst_cellmath__24_0_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_sin_inst_cellmath__66_0_bdw1946085813_bdw cynw_cm_float_sin_I12 (.inst_cellmath__66_0_out0(inst_cellmath__66), .inst_cellmath__66_0_in0(inst_cellmath__24), .inst_cellmath__66_0_in1(inst_cellmath__19), .inst_cellmath__66_0_in2(a_sign));
cynw_cm_float_sin_inst_cellmath__67_0_bdw1946085813_bdw cynw_cm_float_sin_I13 (.inst_cellmath__67_0_out0(inst_cellmath__67), .inst_cellmath__67_0_in0(inst_cellmath__24), .inst_cellmath__67_0_in1(inst_cellmath__19), .inst_cellmath__67_0_in2(a_sign));
cynw_cm_float_sin_inst_cellmath__68_0_bdw1946085813_bdw cynw_cm_float_sin_I14 (.inst_cellmath__68_0_out0(inst_cellmath__68), .inst_cellmath__68_0_in0(inst_cellmath__67), .inst_cellmath__68_0_in1(inst_cellmath__66));
cynw_cm_float_sin_inst_cellmath__69_0_bdw1946085813_bdw cynw_cm_float_sin_I15 (.inst_cellmath__69_0_out0(inst_cellmath__69), .inst_cellmath__69_0_in0(inst_cellmath__24), .inst_cellmath__69_0_in1(inst_cellmath__19));
cynw_cm_float_sin_inst_cellmath__82_0_bdw1946085813_bdw cynw_cm_float_sin_I16 (.inst_cellmath__82_0_out0(inst_cellmath__82), .inst_cellmath__82_0_in0(inst_cellmath__69), .inst_cellmath__82_0_in1(inst_cellmath__19));
cynw_cm_float_sin_inst_cellmath__17_0_bdw1946085813_bdw cynw_cm_float_sin_I17 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_sin_inst_cellmath__79__46__bdw1946085813_bdw cynw_cm_float_sin_I18 (.inst_cellmath__79__46__out0({N487}), .inst_cellmath__79__46__in0(inst_cellmath__68), .inst_cellmath__79__46__in1(inst_cellmath__17));
cynw_cm_float_sin_inst_cellmath__228__231__bdw1946085813_bdw cynw_cm_float_sin_I19 (.inst_cellmath__228__231__out0({N759}), .inst_cellmath__228__231__in0(inst_cellmath__82), .inst_cellmath__228__231__in1({N487}), .inst_cellmath__228__231__in2(inst_cellmath__68));
cynw_cm_float_sin_inst_cellmath__216__184__bdw1946085813_bdw cynw_cm_float_sin_I20 (.inst_cellmath__216__184__out0({N639}), .inst_cellmath__216__184__in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_sin_inst_cellmath__219_0_bdw1946085813_bdw cynw_cm_float_sin_I21 (.inst_cellmath__219_0_out0(inst_cellmath__219), .inst_cellmath__219_0_in0({inst_cellmath__61[22]}), .inst_cellmath__219_0_in1({inst_cellmath__200[48]}));
cynw_cm_float_sin_inst_cellmath__211__182__bdw1946085813_bdw cynw_cm_float_sin_I22 (.inst_cellmath__211__182__out0({N545, N544, N543, N542, N541}), .inst_cellmath__211__182__in0({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_sin_inst_cellmath__215_0_bdw1946085813_bdw cynw_cm_float_sin_I23 (.inst_cellmath__215_0_out0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__215_0_in0({N545, N544, N543, N542, N541}));
cynw_cm_float_sin_inst_cellmath__220__188__bdw1946085813_bdw cynw_cm_float_sin_I24 (.inst_cellmath__220__188__out0({N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679}), .inst_cellmath__220__188__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}), .inst_cellmath__220__188__in1({inst_cellmath__210[22], inst_cellmath__210[21], inst_cellmath__210[20], inst_cellmath__210[19], inst_cellmath__210[18], inst_cellmath__210[17], inst_cellmath__210[16], inst_cellmath__210[15], inst_cellmath__210[14], inst_cellmath__210[13], inst_cellmath__210[12], inst_cellmath__210[11], inst_cellmath__210[10], inst_cellmath__210[9], inst_cellmath__210[8], inst_cellmath__210[7], inst_cellmath__210[6], inst_cellmath__210[5], inst_cellmath__210[4], inst_cellmath__210[3], inst_cellmath__210[2], inst_cellmath__210[1], inst_cellmath__210[0]}));
cynw_cm_float_sin_inst_cellmath__221__195__bdw1946085813_bdw cynw_cm_float_sin_I25 (.inst_cellmath__221__195__out0({N677, N676, N675, N674, N673, N672, N671}), .inst_cellmath__221__195__in0({inst_cellmath__215[4], inst_cellmath__215[3], inst_cellmath__215[2], inst_cellmath__215[1], inst_cellmath__215[0]}));
cynw_cm_float_sin_inst_cellmath__220_2WWMM_bdw1946085813_bdw cynw_cm_float_sin_I26 (.inst_cellmath__220_2WWMM_out0({N670, N3584, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640}), .inst_cellmath__220_2WWMM_in0({N677, N676, N675, N674, N673, N672, N671}), .inst_cellmath__220_2WWMM_in1({N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679}), .inst_cellmath__220_2WWMM_in2(inst_cellmath__219), .inst_cellmath__220_2WWMM_in3({N639}), .inst_cellmath__220_2WWMM_in4({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}), .inst_cellmath__220_2WWMM_in5({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_sin_inst_cellmath__223__208__bdw1946085813_bdw cynw_cm_float_sin_I27 (.inst_cellmath__223__208__out0({N578}), .inst_cellmath__223__208__in0({N3584, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640}));
cynw_cm_float_sin_inst_cellmath__223__207__bdw1946085813_bdw cynw_cm_float_sin_I28 (.inst_cellmath__223__207__out0({N577}), .inst_cellmath__223__207__in0({N757}), .inst_cellmath__223__207__in1(a_sign));
cynw_cm_float_sin_inst_cellmath__223__199__bdw1946085813_bdw cynw_cm_float_sin_I29 (.inst_cellmath__223__199__out0({N579}), .inst_cellmath__223__199__in0(inst_cellmath__82), .inst_cellmath__223__199__in1({N487}), .inst_cellmath__223__199__in2({N578}), .inst_cellmath__223__199__in3({N577}));
cynw_cm_float_sin_inst_cellmath__223_0_bdw1946085813_bdw cynw_cm_float_sin_I30 (.inst_cellmath__223_0_out0(x[31]), .inst_cellmath__223_0_in0({N579}), .inst_cellmath__223_0_in1({N639}), .inst_cellmath__223_0_in2(a_sign));
cynw_cm_float_sin_inst_cellmath__224__212__bdw1946085813_bdw cynw_cm_float_sin_I31 (.inst_cellmath__224__212__out0({N580}), .inst_cellmath__224__212__in0(inst_cellmath__82), .inst_cellmath__224__212__in1({N487}));
cynw_cm_float_sin_inst_cellmath__228_0_bdw1946085813_bdw cynw_cm_float_sin_I32 (.inst_cellmath__228_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__228_0_in0({N759}), .inst_cellmath__228_0_in1({N580}), .inst_cellmath__228_0_in2({N647, N646, N645, N644, N643, N642, N641, N640}));
cynw_cm_float_sin_inst_cellmath__231_0_bdw1946085813_bdw cynw_cm_float_sin_I33 (.inst_cellmath__231_0_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__231_0_in0(inst_cellmath__82), .inst_cellmath__231_0_in1({N759}), .inst_cellmath__231_0_in2({N670, N3584, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648}), .inst_cellmath__231_0_in3({inst_cellmath__210[21]}));
assign inst_cellmath__42[6] = 1'B0;
assign inst_cellmath__42[7] = 1'B0;
assign inst_cellmath__42[8] = 1'B0;
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__200[25] = inst_cellmath__210[0];
assign inst_cellmath__200[26] = inst_cellmath__210[1];
assign inst_cellmath__200[27] = inst_cellmath__210[2];
assign inst_cellmath__200[28] = inst_cellmath__210[3];
assign inst_cellmath__200[29] = inst_cellmath__210[4];
assign inst_cellmath__200[30] = inst_cellmath__210[5];
assign inst_cellmath__200[31] = inst_cellmath__210[6];
assign inst_cellmath__200[32] = inst_cellmath__210[7];
assign inst_cellmath__200[33] = inst_cellmath__210[8];
assign inst_cellmath__200[34] = inst_cellmath__210[9];
assign inst_cellmath__200[35] = inst_cellmath__210[10];
assign inst_cellmath__200[36] = inst_cellmath__210[11];
assign inst_cellmath__200[37] = inst_cellmath__210[12];
assign inst_cellmath__200[38] = inst_cellmath__210[13];
assign inst_cellmath__200[39] = inst_cellmath__210[14];
assign inst_cellmath__200[40] = inst_cellmath__210[15];
assign inst_cellmath__200[41] = inst_cellmath__210[16];
assign inst_cellmath__200[42] = inst_cellmath__210[17];
assign inst_cellmath__200[43] = inst_cellmath__210[18];
assign inst_cellmath__200[44] = inst_cellmath__210[19];
assign inst_cellmath__200[45] = inst_cellmath__210[20];
assign inst_cellmath__200[46] = inst_cellmath__210[21];
assign inst_cellmath__200[47] = inst_cellmath__210[22];
assign inst_cellmath__200[49] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

module cynw_cm_float_sin_inst_blk01_cellmath__39_bdw1946085813_bdw (
	inst_blk01_cellmath__39_out0,
	inst_blk01_cellmath__39_in0
	); /* architecture "gate_level" */ 
output [55:0] inst_blk01_cellmath__39_out0;
input [22:0] inst_blk01_cellmath__39_in0;
wire N354,N360,N362,N366,N368,N370,N372 
	,N374,N376,N378,N380,N382,N384,N386,N388 
	,N390,N392,N394,N396,N1066,N1067,N1070,N1071 
	,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079 
	,N1082,N1083,N1084,N1085,N1088,N1089,N1090,N1091 
	,N1094,N1095,N1096,N1097,N1098,N1099,N1102,N1103 
	,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111 
	,N1114,N1115,N1116,N1117,N1118,N1119,N1122,N1123 
	,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131 
	,N1132,N1133,N1136,N1137,N1138,N1139,N1140,N1141 
	,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149 
	,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157 
	,N1158,N1159,N1160,N1161,N1162,N1163,N1166,N1167 
	,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177 
	,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185 
	,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193 
	,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201 
	,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209 
	,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217 
	,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225 
	,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233 
	,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241 
	,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249 
	,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257 
	,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265 
	,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273 
	,N1274,N1275,N1278,N1279,N1282,N1283,N1286,N1287 
	,N1294,N1295,N1298,N1299,N1300,N1301,N1302,N1303 
	,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311 
	,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319 
	,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327 
	,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335 
	,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343 
	,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351 
	,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359 
	,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367 
	,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375 
	,N1376,N1377,N1378,N1379,N1380,N1381,N1384,N1385 
	,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393 
	,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401 
	,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409 
	,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417 
	,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425 
	,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433 
	,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441 
	,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449 
	,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457 
	,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465 
	,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473 
	,N1474,N1475,N1476,N1477,N1482,N1483,N1484,N1485 
	,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493 
	,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501 
	,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1511 
	,N1521,N1531,N1535,N1536,N1547,N1561,N1565,N1566 
	,N1583,N1611,N1613,N1617,N1618,N1621,N1622,N1661 
	,N1663,N1665,N1684,N1687,N1690,N1693,N1696,N1699 
	,N1702,N1705,N1708,N1711,N1714,N1717,N1734,N1736 
	,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744 
	,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752 
	,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760 
	,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768 
	,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776 
	,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784 
	,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792 
	,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800 
	,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808 
	,N1809,N1810,N1811,N1814,N1818,N1819,N1826,N1830 
	,N1831,N1834,N1835,N1842,N1843,N1846,N1847,N1850 
	,N1851,N1858,N1859,N1862,N1863,N1866,N1867,N1874 
	,N1875,N1878,N1879,N1882,N1883,N1890,N1891,N1894 
	,N1895,N1898,N1899,N1906,N1907,N1910,N1911,N1914 
	,N1915,N1922,N1923,N1926,N1927,N1930,N1931,N1938 
	,N1939,N1942,N1943,N1946,N1947,N1952,N1953,N1954 
	,N1955,N1964,N1966,N1968,N1974,N1975,N2002,N2004 
	,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012 
	,N2013,N2014,N2015,N2020,N2022,N2024,N2025,N2026 
	,N2027,N2028,N2029,N2030,N2031,N2040,N2042,N2044 
	,N2046,N2154,N2157,N2160,N2163,N2166,N2175,N2178 
	,N2187,N2190,N2199,N2202,N2211,N2214,N2223,N2226 
	,N2235,N2238,N2259,N2262,N2278,N2279,N2281,N2282 
	,N2284,N2285,N2287,N2288,N2290,N2291,N2293,N2294 
	,N2296,N2297,N2299,N2300,N2302,N2303,N2305,N2306 
	,N2308,N2309,N2311,N2312,N2314,N2315,N2317,N2318 
	,N2320,N2321,N2323,N2324,N2326,N2327,N2329,N2330 
	,N2332,N2333,N2335,N2336,N2338,N2339,N2341,N2342 
	,N2344,N2345,N2347,N2348,N2350,N2351,N2353,N2354 
	,N2356,N2357,N2553,N2555,N2564,N2566,N2582,N2584 
	,N2593,N2595,N2611,N2613,N2622,N2624,N2640,N2642 
	,N2651,N2653,N2669,N2671,N2680,N2682,N2698,N2700 
	,N2709,N2711,N2727,N2729,N2738,N2740,N2749,N2751 
	,N2760,N2762,N2771,N2773,N2782,N2784,N2800,N2802 
	,N2974,N3013,N3014,N3019,N3022,N3031,N3036,N3037 
	,N3040,N3042,N3043,N3055,N3065,N3073,N3083,N3093 
	,N3101,N3109,N3116,N3117,N3120,N3121,N3133,N3152 
	,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160 
	,N3165,N3170,N3176,N3182,N3188,N3194,N3200,N3206 
	,N3208,N3220,N3221,N3224,N3231,N3238,N3245,N3252 
	,N3259,N3271,N3278,N3285,N3292,N3299,N3306;
INVX2 inst_blk01_cellmath__39_I5 (.Y(N1482), .A(inst_blk01_cellmath__39_in0[0]));
CLKINVX6 inst_blk01_cellmath__39_I6 (.Y(N354), .A(inst_blk01_cellmath__39_in0[1]));
CLKINVX4 inst_blk01_cellmath__39_I7 (.Y(N1484), .A(inst_blk01_cellmath__39_in0[2]));
CLKINVX4 inst_blk01_cellmath__39_I8 (.Y(N1381), .A(inst_blk01_cellmath__39_in0[3]));
CLKINVX6 inst_blk01_cellmath__39_I9 (.Y(N360), .A(inst_blk01_cellmath__39_in0[4]));
CLKINVX6 inst_blk01_cellmath__39_I10 (.Y(N362), .A(inst_blk01_cellmath__39_in0[5]));
CLKINVX12 inst_blk01_cellmath__39_I11 (.Y(N1295), .A(inst_blk01_cellmath__39_in0[6]));
CLKINVX6 inst_blk01_cellmath__39_I12 (.Y(N366), .A(inst_blk01_cellmath__39_in0[7]));
CLKINVX4 inst_blk01_cellmath__39_I13 (.Y(N368), .A(inst_blk01_cellmath__39_in0[8]));
CLKINVX6 inst_blk01_cellmath__39_I14 (.Y(N370), .A(inst_blk01_cellmath__39_in0[9]));
CLKINVX8 inst_blk01_cellmath__39_I15 (.Y(N372), .A(inst_blk01_cellmath__39_in0[10]));
INVX2 inst_blk01_cellmath__39_I16 (.Y(N374), .A(inst_blk01_cellmath__39_in0[11]));
INVX2 inst_blk01_cellmath__39_I17 (.Y(N376), .A(inst_blk01_cellmath__39_in0[12]));
CLKINVX4 inst_blk01_cellmath__39_I18 (.Y(N378), .A(inst_blk01_cellmath__39_in0[13]));
INVX3 inst_blk01_cellmath__39_I19 (.Y(N380), .A(inst_blk01_cellmath__39_in0[14]));
INVX2 inst_blk01_cellmath__39_I20 (.Y(N382), .A(inst_blk01_cellmath__39_in0[15]));
INVX2 inst_blk01_cellmath__39_I21 (.Y(N384), .A(inst_blk01_cellmath__39_in0[16]));
INVX2 inst_blk01_cellmath__39_I22 (.Y(N386), .A(inst_blk01_cellmath__39_in0[17]));
INVX2 inst_blk01_cellmath__39_I23 (.Y(N388), .A(inst_blk01_cellmath__39_in0[18]));
INVX2 inst_blk01_cellmath__39_I24 (.Y(N390), .A(inst_blk01_cellmath__39_in0[19]));
INVX2 inst_blk01_cellmath__39_I25 (.Y(N392), .A(inst_blk01_cellmath__39_in0[20]));
INVX2 inst_blk01_cellmath__39_I26 (.Y(N394), .A(inst_blk01_cellmath__39_in0[21]));
INVXL inst_blk01_cellmath__39_I27 (.Y(N396), .A(inst_blk01_cellmath__39_in0[22]));
BUFX2 inst_blk01_cellmath__39_I1799 (.Y(N2974), .A(N396));
XNOR2X1 hap1_A_I1398 (.Y(N1066), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[2]));
OR2XL hap1_A_I1399 (.Y(N1067), .A(inst_blk01_cellmath__39_in0[9]), .B(inst_blk01_cellmath__39_in0[2]));
ADDFX1 inst_blk01_cellmath__39_I332 (.CO(N1071), .S(N1070), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[10]), .CI(N354));
ADDFHXL inst_blk01_cellmath__39_I333 (.CO(N1073), .S(N1072), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[11]), .CI(N1484));
ADDFXL inst_blk01_cellmath__39_I334 (.CO(N1075), .S(N1074), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[12]), .CI(N1381));
ADDFX1 inst_blk01_cellmath__39_I335 (.CO(N1077), .S(N1076), .A(inst_blk01_cellmath__39_in0[6]), .B(inst_blk01_cellmath__39_in0[13]), .CI(N360));
XNOR2X1 hap1_A_I1400 (.Y(N1078), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[7]));
OR2XL hap1_A_I1401 (.Y(N1079), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[7]));
ADDHX1 inst_blk01_cellmath__39_I337 (.CO(N1083), .S(N1082), .A(N1482), .B(N362));
XNOR2X1 hap1_A_I1402 (.Y(N1084), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[8]));
OR2XL hap1_A_I1403 (.Y(N1085), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[8]));
ADDFHXL inst_blk01_cellmath__39_I339 (.CO(N1089), .S(N1088), .A(N1295), .B(N372), .CI(N354));
XNOR2X1 hap1_A_I1404 (.Y(N1090), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[9]));
OR2XL hap1_A_I1405 (.Y(N1091), .A(inst_blk01_cellmath__39_in0[16]), .B(inst_blk01_cellmath__39_in0[9]));
ADDFX1 inst_blk01_cellmath__39_I341 (.CO(N1095), .S(N1094), .A(N1484), .B(inst_blk01_cellmath__39_in0[0]), .CI(N366));
ADDHX1 inst_blk01_cellmath__39_I342 (.CO(N1097), .S(N1096), .A(N374), .B(N396));
XNOR2X1 hap1_A_I1406 (.Y(N1098), .A(inst_blk01_cellmath__39_in0[17]), .B(inst_blk01_cellmath__39_in0[10]));
OR2XL hap1_A_I1407 (.Y(N1099), .A(inst_blk01_cellmath__39_in0[17]), .B(inst_blk01_cellmath__39_in0[10]));
ADDFX1 inst_blk01_cellmath__39_I344 (.CO(N1103), .S(N1102), .A(N1381), .B(inst_blk01_cellmath__39_in0[1]), .CI(N368));
ADDHX1 inst_blk01_cellmath__39_I345 (.CO(N1105), .S(N1104), .A(N376), .B(N392));
ADDFX1 inst_blk01_cellmath__39_I346 (.CO(N1107), .S(N1106), .A(inst_blk01_cellmath__39_in0[11]), .B(inst_blk01_cellmath__39_in0[18]), .CI(inst_blk01_cellmath__39_in0[2]));
ADDFX1 inst_blk01_cellmath__39_I347 (.CO(N1109), .S(N1108), .A(N370), .B(N360), .CI(N378));
XNOR2X1 hap1_A_I1408 (.Y(N1110), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[12]));
OR2XL hap1_A_I1409 (.Y(N1111), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[12]));
ADDFHXL inst_blk01_cellmath__39_I349 (.CO(N1115), .S(N1114), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[0]), .CI(N362));
ADDHX1 inst_blk01_cellmath__39_I350 (.CO(N1117), .S(N1116), .A(N372), .B(N380));
XNOR2X1 hap1_A_I1410 (.Y(N1118), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[13]));
OR2XL hap1_A_I1411 (.Y(N1119), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[13]));
ADDFX1 inst_blk01_cellmath__39_I352 (.CO(N1123), .S(N1122), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[1]), .CI(N1295));
ADDHX1 inst_blk01_cellmath__39_I353 (.CO(N1125), .S(N1124), .A(N374), .B(N382));
ADDFX1 inst_blk01_cellmath__39_I354 (.CO(N1127), .S(N1126), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[21]), .CI(inst_blk01_cellmath__39_in0[0]));
ADDFHXL inst_blk01_cellmath__39_I355 (.CO(N1129), .S(N1128), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[2]), .CI(N366));
ADDHX1 inst_blk01_cellmath__39_I356 (.CO(N1131), .S(N1130), .A(N376), .B(N384));
XNOR2X1 hap1_A_I1412 (.Y(N1132), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[15]));
OR2XL hap1_A_I1413 (.Y(N1133), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[15]));
ADDFX1 inst_blk01_cellmath__39_I358 (.CO(N1137), .S(N1136), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[1]), .CI(inst_blk01_cellmath__39_in0[6]));
ADDFX1 inst_blk01_cellmath__39_I359 (.CO(N1139), .S(N1138), .A(N378), .B(N368), .CI(N386));
ADDFX1 inst_blk01_cellmath__39_I360 (.CO(N1141), .S(N1140), .A(inst_blk01_cellmath__39_in0[2]), .B(inst_blk01_cellmath__39_in0[16]), .CI(inst_blk01_cellmath__39_in0[4]));
ADDFX1 inst_blk01_cellmath__39_I361 (.CO(N1143), .S(N1142), .A(N370), .B(inst_blk01_cellmath__39_in0[7]), .CI(N380));
ADDFX1 inst_blk01_cellmath__39_I362 (.CO(N1145), .S(N1144), .A(inst_blk01_cellmath__39_in0[3]), .B(inst_blk01_cellmath__39_in0[17]), .CI(inst_blk01_cellmath__39_in0[5]));
ADDHX1 inst_blk01_cellmath__39_I363 (.CO(N1147), .S(N1146), .A(inst_blk01_cellmath__39_in0[8]), .B(N372));
ADDFX1 inst_blk01_cellmath__39_I364 (.CO(N1149), .S(N1148), .A(inst_blk01_cellmath__39_in0[4]), .B(inst_blk01_cellmath__39_in0[18]), .CI(inst_blk01_cellmath__39_in0[6]));
ADDHX1 inst_blk01_cellmath__39_I365 (.CO(N1151), .S(N1150), .A(inst_blk01_cellmath__39_in0[9]), .B(N374));
ADDFX1 inst_blk01_cellmath__39_I366 (.CO(N1153), .S(N1152), .A(inst_blk01_cellmath__39_in0[5]), .B(inst_blk01_cellmath__39_in0[19]), .CI(inst_blk01_cellmath__39_in0[7]));
ADDHX1 inst_blk01_cellmath__39_I367 (.CO(N1155), .S(N1154), .A(inst_blk01_cellmath__39_in0[10]), .B(N376));
ADDFX1 inst_blk01_cellmath__39_I368 (.CO(N1157), .S(N1156), .A(inst_blk01_cellmath__39_in0[6]), .B(inst_blk01_cellmath__39_in0[20]), .CI(inst_blk01_cellmath__39_in0[8]));
ADDHX1 inst_blk01_cellmath__39_I369 (.CO(N1159), .S(N1158), .A(inst_blk01_cellmath__39_in0[11]), .B(N378));
ADDFX1 inst_blk01_cellmath__39_I370 (.CO(N1161), .S(N1160), .A(inst_blk01_cellmath__39_in0[7]), .B(inst_blk01_cellmath__39_in0[21]), .CI(inst_blk01_cellmath__39_in0[9]));
XNOR2X1 hap1_A_I1414 (.Y(N1162), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[8]));
OR2XL hap1_A_I1415 (.Y(N1163), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[8]));
XNOR2X1 hap1_A_I1416 (.Y(N1166), .A(inst_blk01_cellmath__39_in0[5]), .B(N1482));
OR2XL hap1_A_I1417 (.Y(N1167), .A(inst_blk01_cellmath__39_in0[5]), .B(N1482));
ADDFX1 inst_blk01_cellmath__39_I373 (.CO(N1171), .S(N1170), .A(N354), .B(inst_blk01_cellmath__39_in0[6]), .CI(N382));
ADDFX1 inst_blk01_cellmath__39_I374 (.CO(N1173), .S(N1172), .A(inst_blk01_cellmath__39_in0[0]), .B(inst_blk01_cellmath__39_in0[7]), .CI(N1484));
ADDHX1 inst_blk01_cellmath__39_I375 (.CO(N1175), .S(N1174), .A(N384), .B(N378));
ADDFX1 inst_blk01_cellmath__39_I376 (.CO(N1177), .S(N1176), .A(inst_blk01_cellmath__39_in0[1]), .B(inst_blk01_cellmath__39_in0[8]), .CI(N1381));
ADDFX1 inst_blk01_cellmath__39_I377 (.CO(N1179), .S(N1178), .A(N380), .B(N386), .CI(N374));
ADDFX1 inst_blk01_cellmath__39_I378 (.CO(N1181), .S(N1180), .A(N360), .B(N1482), .CI(N388));
ADDFX1 inst_blk01_cellmath__39_I379 (.CO(N1183), .S(N1182), .A(N376), .B(N382), .CI(N1066));
ADDFX1 inst_blk01_cellmath__39_I380 (.CO(N1185), .S(N1184), .A(N384), .B(N362), .CI(N390));
ADDFX1 inst_blk01_cellmath__39_I381 (.CO(N1187), .S(N1186), .A(N1067), .B(N378), .CI(N1070));
ADDFX1 inst_blk01_cellmath__39_I382 (.CO(N1189), .S(N1188), .A(N386), .B(N1295), .CI(N392));
ADDFX1 inst_blk01_cellmath__39_I383 (.CO(N1191), .S(N1190), .A(N1071), .B(N380), .CI(N1072));
ADDFX1 inst_blk01_cellmath__39_I384 (.CO(N1193), .S(N1192), .A(N388), .B(N366), .CI(N394));
ADDFX1 inst_blk01_cellmath__39_I385 (.CO(N1195), .S(N1194), .A(N1073), .B(N382), .CI(N1074));
ADDFXL inst_blk01_cellmath__39_I386 (.CO(N1197), .S(N1196), .A(N2974), .B(N368), .CI(N390));
ADDFHXL inst_blk01_cellmath__39_I387 (.CO(N1199), .S(N1198), .A(N1075), .B(N384), .CI(N1076));
ADDFX1 inst_blk01_cellmath__39_I388 (.CO(N1201), .S(N1200), .A(N392), .B(N370), .CI(N386));
ADDFX1 inst_blk01_cellmath__39_I389 (.CO(N1203), .S(N1202), .A(N1082), .B(N1077), .CI(N1078));
ADDFX1 inst_blk01_cellmath__39_I390 (.CO(N1205), .S(N1204), .A(N388), .B(N394), .CI(N1079));
ADDFX1 inst_blk01_cellmath__39_I391 (.CO(N1207), .S(N1206), .A(N1084), .B(N1083), .CI(N1088));
ADDFHXL inst_blk01_cellmath__39_I392 (.CO(N1209), .S(N1208), .A(N1085), .B(N390), .CI(N1089));
ADDFX1 inst_blk01_cellmath__39_I393 (.CO(N1211), .S(N1210), .A(N1090), .B(N1096), .CI(N1094));
ADDFX1 inst_blk01_cellmath__39_I394 (.CO(N1213), .S(N1212), .A(N1097), .B(N1091), .CI(N1095));
ADDFXL inst_blk01_cellmath__39_I395 (.CO(N1215), .S(N1214), .A(N1098), .B(N1104), .CI(N1102));
ADDFX1 inst_blk01_cellmath__39_I396 (.CO(N1217), .S(N1216), .A(N1099), .B(N394), .CI(N1105));
ADDFX1 inst_blk01_cellmath__39_I397 (.CO(N1219), .S(N1218), .A(N1106), .B(N1103), .CI(N1108));
ADDFXL inst_blk01_cellmath__39_I398 (.CO(N1221), .S(N1220), .A(N1107), .B(N2974), .CI(N1109));
ADDFX1 inst_blk01_cellmath__39_I399 (.CO(N1223), .S(N1222), .A(N1116), .B(N1110), .CI(N1114));
ADDFX1 inst_blk01_cellmath__39_I400 (.CO(N1225), .S(N1224), .A(N1117), .B(N1111), .CI(N1115));
ADDFX1 inst_blk01_cellmath__39_I401 (.CO(N1227), .S(N1226), .A(N1118), .B(N1124), .CI(N1122));
ADDFX1 inst_blk01_cellmath__39_I402 (.CO(N1229), .S(N1228), .A(N1125), .B(N1119), .CI(N1123));
ADDFX1 inst_blk01_cellmath__39_I403 (.CO(N1231), .S(N1230), .A(N1126), .B(N1128), .CI(N1130));
ADDFXL inst_blk01_cellmath__39_I404 (.CO(N1233), .S(N1232), .A(N1129), .B(N1127), .CI(N1131));
ADDFX1 inst_blk01_cellmath__39_I405 (.CO(N1235), .S(N1234), .A(N1136), .B(N1132), .CI(N1138));
ADDFX1 inst_blk01_cellmath__39_I406 (.CO(N1237), .S(N1236), .A(N1133), .B(N388), .CI(N1137));
ADDFXL inst_blk01_cellmath__39_I407 (.CO(N1239), .S(N1238), .A(N1140), .B(N1139), .CI(N1142));
ADDFX1 inst_blk01_cellmath__39_I408 (.CO(N1241), .S(N1240), .A(N390), .B(N382), .CI(N1141));
ADDFX1 inst_blk01_cellmath__39_I409 (.CO(N1243), .S(N1242), .A(N1143), .B(N1146), .CI(N1144));
ADDFX1 inst_blk01_cellmath__39_I410 (.CO(N1245), .S(N1244), .A(N392), .B(N384), .CI(N1147));
ADDFX1 inst_blk01_cellmath__39_I411 (.CO(N1247), .S(N1246), .A(N1150), .B(N1145), .CI(N1148));
ADDFX1 inst_blk01_cellmath__39_I412 (.CO(N1249), .S(N1248), .A(N394), .B(N386), .CI(N1151));
ADDFX1 inst_blk01_cellmath__39_I413 (.CO(N1251), .S(N1250), .A(N1154), .B(N1149), .CI(N1152));
ADDFX1 inst_blk01_cellmath__39_I414 (.CO(N1253), .S(N1252), .A(N2974), .B(N388), .CI(N1155));
ADDFX1 inst_blk01_cellmath__39_I415 (.CO(N1255), .S(N1254), .A(N1158), .B(N1153), .CI(N1156));
ADDFX1 inst_blk01_cellmath__39_I416 (.CO(N1257), .S(N1256), .A(N390), .B(inst_blk01_cellmath__39_in0[12]), .CI(N380));
ADDFX1 inst_blk01_cellmath__39_I417 (.CO(N1259), .S(N1258), .A(N1157), .B(N1159), .CI(N1160));
ADDFX1 inst_blk01_cellmath__39_I418 (.CO(N1261), .S(N1260), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[10]), .CI(N382));
ADDFX1 inst_blk01_cellmath__39_I419 (.CO(N1263), .S(N1262), .A(N1161), .B(N392), .CI(N1162));
ADDFX1 inst_blk01_cellmath__39_I420 (.CO(N1265), .S(N1264), .A(inst_blk01_cellmath__39_in0[11]), .B(inst_blk01_cellmath__39_in0[9]), .CI(inst_blk01_cellmath__39_in0[14]));
ADDFX1 inst_blk01_cellmath__39_I421 (.CO(N1267), .S(N1266), .A(N394), .B(N384), .CI(N1163));
ADDFX1 inst_blk01_cellmath__39_I422 (.CO(N1269), .S(N1268), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[10]), .CI(inst_blk01_cellmath__39_in0[15]));
ADDHX1 inst_blk01_cellmath__39_I423 (.CO(N1271), .S(N1270), .A(N386), .B(N2974));
ADDFX1 inst_blk01_cellmath__39_I424 (.CO(N1273), .S(N1272), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[11]), .CI(inst_blk01_cellmath__39_in0[16]));
XNOR2X1 hap1_A_I1418 (.Y(N1274), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[14]));
OR2XL hap1_A_I1419 (.Y(N1275), .A(inst_blk01_cellmath__39_in0[12]), .B(inst_blk01_cellmath__39_in0[14]));
XNOR2X1 hap1_A_I1420 (.Y(N1278), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[15]));
OR2XL hap1_A_I1421 (.Y(N1279), .A(inst_blk01_cellmath__39_in0[13]), .B(inst_blk01_cellmath__39_in0[15]));
XNOR2X1 hap1_A_I1422 (.Y(N1282), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[16]));
OR2XL hap1_A_I1423 (.Y(N1283), .A(inst_blk01_cellmath__39_in0[14]), .B(inst_blk01_cellmath__39_in0[16]));
XNOR2X1 hap1_A_I1424 (.Y(N1286), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[17]));
OR2XL hap1_A_I1425 (.Y(N1287), .A(inst_blk01_cellmath__39_in0[15]), .B(inst_blk01_cellmath__39_in0[17]));
INVXL inst_blk01_cellmath__39_I430 (.Y(N1294), .A(N1295));
ADDHX1 inst_blk01_cellmath__39_I431 (.CO(N1299), .S(N1298), .A(N366), .B(N360));
ADDHX1 inst_blk01_cellmath__39_I432 (.CO(N1301), .S(N1300), .A(N368), .B(N362));
ADDFX1 inst_blk01_cellmath__39_I433 (.CO(N1303), .S(N1302), .A(N370), .B(inst_blk01_cellmath__39_in0[0]), .CI(N1295));
ADDFX1 inst_blk01_cellmath__39_I434 (.CO(N1305), .S(N1304), .A(N372), .B(inst_blk01_cellmath__39_in0[1]), .CI(N366));
ADDFX1 inst_blk01_cellmath__39_I435 (.CO(N1307), .S(N1306), .A(N374), .B(inst_blk01_cellmath__39_in0[2]), .CI(N368));
ADDFX1 inst_blk01_cellmath__39_I436 (.CO(N1309), .S(N1308), .A(N376), .B(inst_blk01_cellmath__39_in0[3]), .CI(N370));
ADDFX1 inst_blk01_cellmath__39_I437 (.CO(N1311), .S(N1310), .A(N378), .B(inst_blk01_cellmath__39_in0[4]), .CI(N372));
ADDFX1 inst_blk01_cellmath__39_I438 (.CO(N1313), .S(N1312), .A(N374), .B(N380), .CI(N368));
ADDFX1 inst_blk01_cellmath__39_I439 (.CO(N1315), .S(N1314), .A(N370), .B(N376), .CI(N1167));
ADDFX1 inst_blk01_cellmath__39_I440 (.CO(N1317), .S(N1316), .A(N1174), .B(N372), .CI(N1171));
ADDFX1 inst_blk01_cellmath__39_I441 (.CO(N1319), .S(N1318), .A(N1173), .B(N1175), .CI(N1176));
ADDFX1 inst_blk01_cellmath__39_I442 (.CO(N1321), .S(N1320), .A(N1179), .B(N1177), .CI(N1180));
ADDFX1 inst_blk01_cellmath__39_I443 (.CO(N1323), .S(N1322), .A(N1184), .B(N1181), .CI(N1183));
ADDFX1 inst_blk01_cellmath__39_I444 (.CO(N1325), .S(N1324), .A(N1188), .B(N1185), .CI(N1187));
ADDFHXL inst_blk01_cellmath__39_I445 (.CO(N1327), .S(N1326), .A(N1192), .B(N1189), .CI(N1191));
ADDFXL inst_blk01_cellmath__39_I446 (.CO(N1329), .S(N1328), .A(N1196), .B(N1193), .CI(N1195));
ADDFHXL inst_blk01_cellmath__39_I447 (.CO(N1331), .S(N1330), .A(N1200), .B(N1197), .CI(N1199));
ADDFX1 inst_blk01_cellmath__39_I448 (.CO(N1333), .S(N1332), .A(N1204), .B(N1201), .CI(N1203));
ADDFHXL inst_blk01_cellmath__39_I449 (.CO(N1335), .S(N1334), .A(N1208), .B(N1205), .CI(N1207));
ADDFXL inst_blk01_cellmath__39_I450 (.CO(N1337), .S(N1336), .A(N1212), .B(N1209), .CI(N1211));
ADDFHXL inst_blk01_cellmath__39_I451 (.CO(N1339), .S(N1338), .A(N1216), .B(N1213), .CI(N1215));
ADDFHXL inst_blk01_cellmath__39_I452 (.CO(N1341), .S(N1340), .A(N1220), .B(N1217), .CI(N1219));
ADDFXL inst_blk01_cellmath__39_I453 (.CO(N1343), .S(N1342), .A(N1223), .B(N1221), .CI(N1224));
ADDFXL inst_blk01_cellmath__39_I454 (.CO(N1345), .S(N1344), .A(N1227), .B(N1225), .CI(N1228));
ADDFXL inst_blk01_cellmath__39_I455 (.CO(N1347), .S(N1346), .A(N1232), .B(N1229), .CI(N1231));
ADDFHXL inst_blk01_cellmath__39_I456 (.CO(N1349), .S(N1348), .A(N1236), .B(N1233), .CI(N1235));
ADDFHXL inst_blk01_cellmath__39_I457 (.CO(N1351), .S(N1350), .A(N1240), .B(N1237), .CI(N1239));
ADDFX1 inst_blk01_cellmath__39_I458 (.CO(N1353), .S(N1352), .A(N1244), .B(N1241), .CI(N1243));
ADDFX1 inst_blk01_cellmath__39_I459 (.CO(N1355), .S(N1354), .A(N1248), .B(N1245), .CI(N1247));
ADDFX1 inst_blk01_cellmath__39_I460 (.CO(N1357), .S(N1356), .A(N1252), .B(N1249), .CI(N1251));
ADDFXL inst_blk01_cellmath__39_I461 (.CO(N1359), .S(N1358), .A(N1253), .B(N1256), .CI(N1255));
ADDFX1 inst_blk01_cellmath__39_I462 (.CO(N1361), .S(N1360), .A(N1260), .B(N1257), .CI(N1259));
ADDFX1 inst_blk01_cellmath__39_I463 (.CO(N1363), .S(N1362), .A(N1264), .B(N1261), .CI(N1263));
ADDFX1 inst_blk01_cellmath__39_I464 (.CO(N1365), .S(N1364), .A(N1270), .B(N1265), .CI(N1268));
ADDFX1 inst_blk01_cellmath__39_I465 (.CO(N1367), .S(N1366), .A(N1271), .B(N388), .CI(N1269));
ADDFX1 inst_blk01_cellmath__39_I466 (.CO(N1369), .S(N1368), .A(N390), .B(inst_blk01_cellmath__39_in0[17]), .CI(N1273));
ADDFX1 inst_blk01_cellmath__39_I467 (.CO(N1371), .S(N1370), .A(N392), .B(inst_blk01_cellmath__39_in0[18]), .CI(N1275));
ADDFX1 inst_blk01_cellmath__39_I468 (.CO(N1373), .S(N1372), .A(N394), .B(inst_blk01_cellmath__39_in0[19]), .CI(N1279));
ADDFX1 inst_blk01_cellmath__39_I469 (.CO(N1375), .S(N1374), .A(N2974), .B(inst_blk01_cellmath__39_in0[20]), .CI(N1283));
ADDFX1 inst_blk01_cellmath__39_I470 (.CO(N1377), .S(N1376), .A(inst_blk01_cellmath__39_in0[21]), .B(inst_blk01_cellmath__39_in0[18]), .CI(N384));
ADDFX1 inst_blk01_cellmath__39_I471 (.CO(N1379), .S(N1378), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[17]), .CI(inst_blk01_cellmath__39_in0[22]));
INVXL inst_blk01_cellmath__39_I472 (.Y(N1380), .A(N1381));
ADDHX1 inst_blk01_cellmath__39_I473 (.CO(N1385), .S(N1384), .A(N360), .B(N354));
ADDHX1 inst_blk01_cellmath__39_I474 (.CO(N1387), .S(N1386), .A(N362), .B(N1484));
ADDFX1 inst_blk01_cellmath__39_I475 (.CO(N1389), .S(N1388), .A(N1482), .B(N1381), .CI(N1294));
ADDFX1 inst_blk01_cellmath__39_I476 (.CO(N1391), .S(N1390), .A(N354), .B(N1295), .CI(N1298));
ADDFX1 inst_blk01_cellmath__39_I477 (.CO(N1393), .S(N1392), .A(N1299), .B(N1484), .CI(N1300));
ADDFX1 inst_blk01_cellmath__39_I478 (.CO(N1395), .S(N1394), .A(N1301), .B(N1381), .CI(N1302));
ADDFX1 inst_blk01_cellmath__39_I479 (.CO(N1397), .S(N1396), .A(N1303), .B(N360), .CI(N1304));
ADDFX1 inst_blk01_cellmath__39_I480 (.CO(N1399), .S(N1398), .A(N1305), .B(N362), .CI(N1306));
ADDFX1 inst_blk01_cellmath__39_I481 (.CO(N1401), .S(N1400), .A(N1307), .B(N1295), .CI(N1308));
ADDFX1 inst_blk01_cellmath__39_I482 (.CO(N1403), .S(N1402), .A(N1309), .B(N366), .CI(N1310));
ADDFX1 inst_blk01_cellmath__39_I483 (.CO(N1405), .S(N1404), .A(N1166), .B(N1311), .CI(N1312));
ADDFX1 inst_blk01_cellmath__39_I484 (.CO(N1407), .S(N1406), .A(N1170), .B(N1313), .CI(N1314));
ADDFX1 inst_blk01_cellmath__39_I485 (.CO(N1409), .S(N1408), .A(N1315), .B(N1172), .CI(N1316));
ADDFX1 inst_blk01_cellmath__39_I486 (.CO(N1411), .S(N1410), .A(N1317), .B(N1178), .CI(N1318));
ADDFX1 inst_blk01_cellmath__39_I487 (.CO(N1413), .S(N1412), .A(N1182), .B(N1319), .CI(N1320));
ADDFX1 inst_blk01_cellmath__39_I488 (.CO(N1415), .S(N1414), .A(N1186), .B(N1321), .CI(N1322));
ADDFHXL inst_blk01_cellmath__39_I489 (.CO(N1417), .S(N1416), .A(N1323), .B(N1190), .CI(N1324));
ADDFX1 inst_blk01_cellmath__39_I490 (.CO(N1419), .S(N1418), .A(N1325), .B(N1194), .CI(N1326));
ADDFX1 inst_blk01_cellmath__39_I491 (.CO(N1421), .S(N1420), .A(N1327), .B(N1198), .CI(N1328));
ADDFHXL inst_blk01_cellmath__39_I492 (.CO(N1423), .S(N1422), .A(N1329), .B(N1202), .CI(N1330));
ADDFX1 inst_blk01_cellmath__39_I493 (.CO(N1425), .S(N1424), .A(N1331), .B(N1206), .CI(N1332));
ADDFHX1 inst_blk01_cellmath__39_I494 (.CO(N1427), .S(N1426), .A(N1333), .B(N1210), .CI(N1334));
ADDFHXL inst_blk01_cellmath__39_I495 (.CO(N1429), .S(N1428), .A(N1335), .B(N1214), .CI(N1336));
ADDFHX1 inst_blk01_cellmath__39_I496 (.CO(N1431), .S(N1430), .A(N1337), .B(N1218), .CI(N1338));
ADDFHX1 inst_blk01_cellmath__39_I497 (.CO(N1433), .S(N1432), .A(N1339), .B(N1222), .CI(N1340));
ADDFHX1 inst_blk01_cellmath__39_I498 (.CO(N1435), .S(N1434), .A(N1341), .B(N1226), .CI(N1342));
ADDFX1 inst_blk01_cellmath__39_I499 (.CO(N1437), .S(N1436), .A(N1343), .B(N1230), .CI(N1344));
ADDFHXL inst_blk01_cellmath__39_I500 (.CO(N1439), .S(N1438), .A(N1345), .B(N1234), .CI(N1346));
ADDFHXL inst_blk01_cellmath__39_I501 (.CO(N1441), .S(N1440), .A(N1347), .B(N1238), .CI(N1348));
ADDFHX1 inst_blk01_cellmath__39_I502 (.CO(N1443), .S(N1442), .A(N1349), .B(N1242), .CI(N1350));
ADDFX1 inst_blk01_cellmath__39_I503 (.CO(N1445), .S(N1444), .A(N1351), .B(N1246), .CI(N1352));
ADDFX1 inst_blk01_cellmath__39_I504 (.CO(N1447), .S(N1446), .A(N1353), .B(N1250), .CI(N1354));
ADDFX1 inst_blk01_cellmath__39_I505 (.CO(N1449), .S(N1448), .A(N1355), .B(N1254), .CI(N1356));
ADDFX1 inst_blk01_cellmath__39_I506 (.CO(N1451), .S(N1450), .A(N1357), .B(N1258), .CI(N1358));
ADDFX1 inst_blk01_cellmath__39_I507 (.CO(N1453), .S(N1452), .A(N1359), .B(N1262), .CI(N1360));
ADDFX1 inst_blk01_cellmath__39_I508 (.CO(N1455), .S(N1454), .A(N1361), .B(N1266), .CI(N1362));
ADDFX1 inst_blk01_cellmath__39_I509 (.CO(N1457), .S(N1456), .A(N1364), .B(N1267), .CI(N1363));
ADDFX1 inst_blk01_cellmath__39_I510 (.CO(N1459), .S(N1458), .A(N1366), .B(N1272), .CI(N1365));
ADDFX1 inst_blk01_cellmath__39_I511 (.CO(N1461), .S(N1460), .A(N1367), .B(N1274), .CI(N1368));
ADDFX1 inst_blk01_cellmath__39_I512 (.CO(N1463), .S(N1462), .A(N1369), .B(N1278), .CI(N1370));
ADDFX1 inst_blk01_cellmath__39_I513 (.CO(N1465), .S(N1464), .A(N1371), .B(N1282), .CI(N1372));
ADDFX1 inst_blk01_cellmath__39_I514 (.CO(N1467), .S(N1466), .A(N1373), .B(N1286), .CI(N1374));
ADDFX1 inst_blk01_cellmath__39_I515 (.CO(N1469), .S(N1468), .A(N1376), .B(N1287), .CI(N1375));
ADDFX1 inst_blk01_cellmath__39_I516 (.CO(N1471), .S(N1470), .A(N1377), .B(inst_blk01_cellmath__39_in0[16]), .CI(N1378));
ADDFX1 inst_blk01_cellmath__39_I517 (.CO(N1473), .S(N1472), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[18]), .CI(N1379));
ADDHX1 inst_blk01_cellmath__39_I518 (.CO(N1475), .S(N1474), .A(inst_blk01_cellmath__39_in0[19]), .B(inst_blk01_cellmath__39_in0[21]));
ADDHX1 inst_blk01_cellmath__39_I519 (.CO(N1477), .S(N1476), .A(inst_blk01_cellmath__39_in0[20]), .B(inst_blk01_cellmath__39_in0[22]));
INVX1 inst_blk01_cellmath__39_I1555 (.Y(inst_blk01_cellmath__39_out0[1]), .A(N1482));
INVXL inst_blk01_cellmath__39_I522 (.Y(N1483), .A(N354));
NOR2XL inst_blk01_cellmath__39_I524 (.Y(N1485), .A(N1482), .B(N1380));
NAND2XL inst_blk01_cellmath__39_I525 (.Y(N1486), .A(N1482), .B(N1380));
NOR2XL inst_blk01_cellmath__39_I526 (.Y(N1487), .A(N1381), .B(N1384));
NAND2XL inst_blk01_cellmath__39_I527 (.Y(N1488), .A(N1381), .B(N1384));
NOR2XL inst_blk01_cellmath__39_I528 (.Y(N1489), .A(N1385), .B(N1386));
NAND2XL inst_blk01_cellmath__39_I529 (.Y(N1490), .A(N1385), .B(N1386));
NOR2XL inst_blk01_cellmath__39_I530 (.Y(N1491), .A(N1387), .B(N1388));
NAND2XL inst_blk01_cellmath__39_I531 (.Y(N1492), .A(N1387), .B(N1388));
NOR2XL inst_blk01_cellmath__39_I532 (.Y(N1493), .A(N1389), .B(N1390));
NAND2XL inst_blk01_cellmath__39_I533 (.Y(N1494), .A(N1389), .B(N1390));
NOR2XL inst_blk01_cellmath__39_I534 (.Y(N1495), .A(N1391), .B(N1392));
NAND2XL inst_blk01_cellmath__39_I535 (.Y(N1496), .A(N1391), .B(N1392));
NOR2XL inst_blk01_cellmath__39_I536 (.Y(N1497), .A(N1393), .B(N1394));
NAND2XL inst_blk01_cellmath__39_I537 (.Y(N1498), .A(N1393), .B(N1394));
NOR2XL inst_blk01_cellmath__39_I538 (.Y(N1499), .A(N1395), .B(N1396));
NAND2XL inst_blk01_cellmath__39_I539 (.Y(N1500), .A(N1395), .B(N1396));
NOR2X1 inst_blk01_cellmath__39_I540 (.Y(N1501), .A(N1397), .B(N1398));
NAND2XL inst_blk01_cellmath__39_I541 (.Y(N1502), .A(N1397), .B(N1398));
NOR2XL inst_blk01_cellmath__39_I542 (.Y(N1503), .A(N1399), .B(N1400));
NAND2X1 inst_blk01_cellmath__39_I543 (.Y(N1504), .A(N1399), .B(N1400));
NOR2XL inst_blk01_cellmath__39_I544 (.Y(N1505), .A(N1401), .B(N1402));
NAND2XL inst_blk01_cellmath__39_I545 (.Y(N1506), .A(N1401), .B(N1402));
NOR2XL inst_blk01_cellmath__39_I546 (.Y(N1507), .A(N1403), .B(N1404));
NAND2XL inst_blk01_cellmath__39_I547 (.Y(N1508), .A(N1403), .B(N1404));
NOR2XL inst_blk01_cellmath__39_I550 (.Y(N1511), .A(N1483), .B(inst_blk01_cellmath__39_out0[1]));
NAND2XL inst_blk01_cellmath__39_I558 (.Y(N1521), .A(N1484), .B(N1511));
AOI21XL inst_blk01_cellmath__39_I566 (.Y(N1531), .A0(N1486), .A1(N1521), .B0(N1485));
AOI21XL inst_blk01_cellmath__39_I570 (.Y(N1535), .A0(N1490), .A1(N1487), .B0(N1489));
NAND2XL inst_blk01_cellmath__39_I571 (.Y(N1536), .A(N1490), .B(N1488));
OAI21XL inst_blk01_cellmath__39_I582 (.Y(N1547), .A0(N1536), .A1(N1531), .B0(N1535));
AOI21XL inst_blk01_cellmath__39_I596 (.Y(N1561), .A0(N1492), .A1(N1547), .B0(N1491));
AOI21XL inst_blk01_cellmath__39_I600 (.Y(N1565), .A0(N1496), .A1(N1493), .B0(N1495));
NAND2XL inst_blk01_cellmath__39_I601 (.Y(N1566), .A(N1496), .B(N1494));
OAI21X1 inst_blk01_cellmath__39_I618 (.Y(N1583), .A0(N1566), .A1(N1561), .B0(N1565));
AO21XL inst_blk01_cellmath__39_I1802 (.Y(N3013), .A0(N1500), .A1(N1497), .B0(N1499));
AND2XL inst_blk01_cellmath__39_I1803 (.Y(N3014), .A(N1500), .B(N1498));
NOR2BX1 andori2bb1_A_I3258 (.Y(N3224), .AN(N1488), .B(N1531));
NOR2XL andori2bb1_A_I1895 (.Y(N3019), .A(N3224), .B(N1487));
NOR2BX1 andori2bb1_A_I3259 (.Y(N3231), .AN(N1494), .B(N1561));
NOR2XL andori2bb1_A_I1897 (.Y(N3022), .A(N3231), .B(N1493));
AOI21XL inst_blk01_cellmath__39_I646 (.Y(N1611), .A0(N1498), .A1(N1583), .B0(N1497));
AOI21X2 inst_blk01_cellmath__39_I648 (.Y(N1613), .A0(N3014), .A1(N1583), .B0(N3013));
AOI21XL inst_blk01_cellmath__39_I652 (.Y(N1617), .A0(N1504), .A1(N1501), .B0(N1503));
NAND2XL inst_blk01_cellmath__39_I653 (.Y(N1618), .A(N1504), .B(N1502));
INVXL inst_blk01_cellmath__39_I1607 (.Y(N3031), .A(N1506));
AOI21XL inst_blk01_cellmath__39_I656 (.Y(N1621), .A0(N1508), .A1(N1505), .B0(N1507));
NAND2XL inst_blk01_cellmath__39_I657 (.Y(N1622), .A(N1508), .B(N1506));
INVXL inst_blk01_cellmath__39_I1612 (.Y(N3036), .A(N1501));
INVXL inst_blk01_cellmath__39_I1613 (.Y(N3037), .A(N1502));
NOR2XL andori2bb1_A_I1898 (.Y(N3238), .A(N3031), .B(N1617));
NOR2XL andori2bb1_A_I1899 (.Y(N3040), .A(N3238), .B(N1505));
OA21X1 inst_blk01_cellmath__39_I1809 (.Y(N3042), .A0(N1622), .A1(N1617), .B0(N1621));
OR2XL inst_blk01_cellmath__39_I1810 (.Y(N3043), .A(N1622), .B(N1618));
OAI21XL inst_blk01_cellmath__39_I696 (.Y(N1661), .A0(N3037), .A1(N1613), .B0(N3036));
OAI21XL inst_blk01_cellmath__39_I698 (.Y(N1663), .A0(N1618), .A1(N1613), .B0(N1617));
OAI31X1 inst_blk01_cellmath__39_I1812 (.Y(N1665), .A0(N3031), .A1(N1618), .A2(N1613), .B0(N3040));
OAI21X1 inst_blk01_cellmath__39_I702 (.Y(N1734), .A0(N3043), .A1(N1613), .B0(N3042));
NAND2BXL inst_blk01_cellmath__39_I715 (.Y(N1684), .AN(N1485), .B(N1486));
NAND2BXL inst_blk01_cellmath__39_I718 (.Y(N1687), .AN(N1487), .B(N1488));
NAND2BXL inst_blk01_cellmath__39_I721 (.Y(N1690), .AN(N1489), .B(N1490));
NAND2BXL inst_blk01_cellmath__39_I724 (.Y(N1693), .AN(N1491), .B(N1492));
NAND2BXL inst_blk01_cellmath__39_I727 (.Y(N1696), .AN(N1493), .B(N1494));
NAND2BXL inst_blk01_cellmath__39_I730 (.Y(N1699), .AN(N1495), .B(N1496));
NAND2BXL inst_blk01_cellmath__39_I733 (.Y(N1702), .AN(N1497), .B(N1498));
NAND2BXL inst_blk01_cellmath__39_I736 (.Y(N1705), .AN(N1499), .B(N1500));
NAND2BXL inst_blk01_cellmath__39_I739 (.Y(N1708), .AN(N1501), .B(N1502));
NAND2BXL inst_blk01_cellmath__39_I742 (.Y(N1711), .AN(N1503), .B(N1504));
NAND2BXL inst_blk01_cellmath__39_I745 (.Y(N1714), .AN(N1505), .B(N1506));
NAND2BXL inst_blk01_cellmath__39_I748 (.Y(N1717), .AN(N1507), .B(N1508));
XOR2XL inst_blk01_cellmath__39_I3262 (.Y(inst_blk01_cellmath__39_out0[2]), .A(inst_blk01_cellmath__39_out0[1]), .B(N1483));
XOR2XL inst_blk01_cellmath__39_I1815 (.Y(inst_blk01_cellmath__39_out0[3]), .A(N1511), .B(N1484));
XOR2XL inst_blk01_cellmath__39_I1816 (.Y(inst_blk01_cellmath__39_out0[4]), .A(N1521), .B(N1684));
XNOR2X1 inst_blk01_cellmath__39_I753 (.Y(inst_blk01_cellmath__39_out0[5]), .A(N1531), .B(N1687));
XNOR2X1 inst_blk01_cellmath__39_I754 (.Y(inst_blk01_cellmath__39_out0[6]), .A(N3019), .B(N1690));
XOR2XL inst_blk01_cellmath__39_I1817 (.Y(inst_blk01_cellmath__39_out0[7]), .A(N1547), .B(N1693));
XNOR2X1 inst_blk01_cellmath__39_I756 (.Y(inst_blk01_cellmath__39_out0[8]), .A(N1561), .B(N1696));
XNOR2X1 inst_blk01_cellmath__39_I757 (.Y(inst_blk01_cellmath__39_out0[9]), .A(N3022), .B(N1699));
XOR2XL inst_blk01_cellmath__39_I1818 (.Y(inst_blk01_cellmath__39_out0[10]), .A(N1583), .B(N1702));
XNOR2X1 inst_blk01_cellmath__39_I759 (.Y(inst_blk01_cellmath__39_out0[11]), .A(N1611), .B(N1705));
XNOR2X1 inst_blk01_cellmath__39_I760 (.Y(inst_blk01_cellmath__39_out0[12]), .A(N1613), .B(N1708));
XOR2XL inst_blk01_cellmath__39_I761 (.Y(inst_blk01_cellmath__39_out0[13]), .A(N1661), .B(N1711));
XOR2XL inst_blk01_cellmath__39_I762 (.Y(inst_blk01_cellmath__39_out0[14]), .A(N1663), .B(N1714));
XOR2XL inst_blk01_cellmath__39_I763 (.Y(inst_blk01_cellmath__39_out0[15]), .A(N1665), .B(N1717));
NOR2XL inst_blk01_cellmath__39_I766 (.Y(N1736), .A(N1405), .B(N1406));
NAND2XL inst_blk01_cellmath__39_I767 (.Y(N1737), .A(N1405), .B(N1406));
NOR2XL inst_blk01_cellmath__39_I768 (.Y(N1738), .A(N1407), .B(N1408));
NAND2XL inst_blk01_cellmath__39_I769 (.Y(N1739), .A(N1407), .B(N1408));
NOR2XL inst_blk01_cellmath__39_I770 (.Y(N1740), .A(N1409), .B(N1410));
NAND2XL inst_blk01_cellmath__39_I771 (.Y(N1741), .A(N1409), .B(N1410));
NOR2X1 inst_blk01_cellmath__39_I772 (.Y(N1742), .A(N1411), .B(N1412));
NAND2XL inst_blk01_cellmath__39_I773 (.Y(N1743), .A(N1411), .B(N1412));
NOR2XL inst_blk01_cellmath__39_I774 (.Y(N1744), .A(N1413), .B(N1414));
NAND2X1 inst_blk01_cellmath__39_I775 (.Y(N1745), .A(N1413), .B(N1414));
NOR2X2 inst_blk01_cellmath__39_I776 (.Y(N1746), .A(N1415), .B(N1416));
NAND2X2 inst_blk01_cellmath__39_I777 (.Y(N1747), .A(N1415), .B(N1416));
NOR2XL inst_blk01_cellmath__39_I778 (.Y(N1748), .A(N1417), .B(N1418));
NAND2X4 inst_blk01_cellmath__39_I779 (.Y(N1749), .A(N1417), .B(N1418));
NOR2X2 inst_blk01_cellmath__39_I780 (.Y(N1750), .A(N1419), .B(N1420));
NAND2X1 inst_blk01_cellmath__39_I781 (.Y(N1751), .A(N1419), .B(N1420));
NOR2X1 inst_blk01_cellmath__39_I782 (.Y(N1752), .A(N1421), .B(N1422));
NAND2X4 inst_blk01_cellmath__39_I783 (.Y(N1753), .A(N1421), .B(N1422));
NOR2X1 inst_blk01_cellmath__39_I784 (.Y(N1754), .A(N1423), .B(N1424));
NAND2X2 inst_blk01_cellmath__39_I785 (.Y(N1755), .A(N1423), .B(N1424));
NOR2X1 inst_blk01_cellmath__39_I1819 (.Y(N1756), .A(N1426), .B(N1425));
NAND2X4 inst_blk01_cellmath__39_I787 (.Y(N1757), .A(N1425), .B(N1426));
NOR2X4 inst_blk01_cellmath__39_I788 (.Y(N1758), .A(N1427), .B(N1428));
NAND2X2 inst_blk01_cellmath__39_I789 (.Y(N1759), .A(N1427), .B(N1428));
NOR2X1 inst_blk01_cellmath__39_I790 (.Y(N1760), .A(N1429), .B(N1430));
NAND2X4 inst_blk01_cellmath__39_I791 (.Y(N1761), .A(N1429), .B(N1430));
NOR2X2 inst_blk01_cellmath__39_I792 (.Y(N1762), .A(N1431), .B(N1432));
NAND2X4 inst_blk01_cellmath__39_I793 (.Y(N1763), .A(N1431), .B(N1432));
NOR2X1 inst_blk01_cellmath__39_I794 (.Y(N1764), .A(N1433), .B(N1434));
NAND2X6 inst_blk01_cellmath__39_I795 (.Y(N1765), .A(N1433), .B(N1434));
NOR2X4 inst_blk01_cellmath__39_I796 (.Y(N1766), .A(N1435), .B(N1436));
NAND2X2 inst_blk01_cellmath__39_I797 (.Y(N1767), .A(N1435), .B(N1436));
NOR2X1 inst_blk01_cellmath__39_I1820 (.Y(N1768), .A(N1438), .B(N1437));
NAND2X4 inst_blk01_cellmath__39_I799 (.Y(N1769), .A(N1437), .B(N1438));
NOR2X2 inst_blk01_cellmath__39_I800 (.Y(N1770), .A(N1439), .B(N1440));
NAND2X2 inst_blk01_cellmath__39_I801 (.Y(N1771), .A(N1439), .B(N1440));
NOR2X1 inst_blk01_cellmath__39_I802 (.Y(N1772), .A(N1441), .B(N1442));
NAND2X6 inst_blk01_cellmath__39_I803 (.Y(N1773), .A(N1441), .B(N1442));
NOR2X2 inst_blk01_cellmath__39_I804 (.Y(N1774), .A(N1443), .B(N1444));
NAND2X2 inst_blk01_cellmath__39_I805 (.Y(N1775), .A(N1443), .B(N1444));
NOR2X1 inst_blk01_cellmath__39_I806 (.Y(N1776), .A(N1445), .B(N1446));
NAND2X4 inst_blk01_cellmath__39_I807 (.Y(N1777), .A(N1445), .B(N1446));
NOR2X1 inst_blk01_cellmath__39_I808 (.Y(N1778), .A(N1447), .B(N1448));
NAND2X2 inst_blk01_cellmath__39_I809 (.Y(N1779), .A(N1447), .B(N1448));
NOR2XL inst_blk01_cellmath__39_I810 (.Y(N1780), .A(N1449), .B(N1450));
NAND2X4 inst_blk01_cellmath__39_I811 (.Y(N1781), .A(N1449), .B(N1450));
NOR2X2 inst_blk01_cellmath__39_I812 (.Y(N1782), .A(N1451), .B(N1452));
NAND2X2 inst_blk01_cellmath__39_I813 (.Y(N1783), .A(N1451), .B(N1452));
NOR2XL inst_blk01_cellmath__39_I814 (.Y(N1784), .A(N1453), .B(N1454));
NAND2X2 inst_blk01_cellmath__39_I815 (.Y(N1785), .A(N1453), .B(N1454));
NOR2XL inst_blk01_cellmath__39_I816 (.Y(N1786), .A(N1455), .B(N1456));
NAND2XL inst_blk01_cellmath__39_I817 (.Y(N1787), .A(N1455), .B(N1456));
NOR2XL inst_blk01_cellmath__39_I818 (.Y(N1788), .A(N1458), .B(N1457));
NAND2X1 inst_blk01_cellmath__39_I819 (.Y(N1789), .A(N1458), .B(N1457));
NOR2XL inst_blk01_cellmath__39_I820 (.Y(N1790), .A(N1459), .B(N1460));
NAND2XL inst_blk01_cellmath__39_I821 (.Y(N1791), .A(N1459), .B(N1460));
NOR2XL inst_blk01_cellmath__39_I822 (.Y(N1792), .A(N1461), .B(N1462));
NAND2XL inst_blk01_cellmath__39_I823 (.Y(N1793), .A(N1461), .B(N1462));
NOR2XL inst_blk01_cellmath__39_I824 (.Y(N1794), .A(N1463), .B(N1464));
NAND2XL inst_blk01_cellmath__39_I825 (.Y(N1795), .A(N1463), .B(N1464));
NOR2XL inst_blk01_cellmath__39_I826 (.Y(N1796), .A(N1465), .B(N1466));
NAND2XL inst_blk01_cellmath__39_I827 (.Y(N1797), .A(N1465), .B(N1466));
NOR2XL inst_blk01_cellmath__39_I828 (.Y(N1798), .A(N1467), .B(N1468));
NAND2XL inst_blk01_cellmath__39_I829 (.Y(N1799), .A(N1467), .B(N1468));
NOR2XL inst_blk01_cellmath__39_I830 (.Y(N1800), .A(N1469), .B(N1470));
NAND2XL inst_blk01_cellmath__39_I831 (.Y(N1801), .A(N1469), .B(N1470));
NOR2XL inst_blk01_cellmath__39_I832 (.Y(N1802), .A(N1472), .B(N1471));
NAND2XL inst_blk01_cellmath__39_I833 (.Y(N1803), .A(N1472), .B(N1471));
NOR2XL inst_blk01_cellmath__39_I834 (.Y(N1804), .A(N1474), .B(N1473));
NAND2XL inst_blk01_cellmath__39_I835 (.Y(N1805), .A(N1474), .B(N1473));
NOR2XL inst_blk01_cellmath__39_I836 (.Y(N1806), .A(N1475), .B(N1476));
NAND2XL inst_blk01_cellmath__39_I837 (.Y(N1807), .A(N1475), .B(N1476));
NOR2XL inst_blk01_cellmath__39_I838 (.Y(N1808), .A(N394), .B(N1477));
NAND2XL inst_blk01_cellmath__39_I839 (.Y(N1809), .A(N394), .B(N1477));
NOR2XL inst_blk01_cellmath__39_I840 (.Y(N1810), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[21]));
NAND2XL inst_blk01_cellmath__39_I841 (.Y(N1811), .A(inst_blk01_cellmath__39_in0[22]), .B(inst_blk01_cellmath__39_in0[21]));
AOI21X1 inst_blk01_cellmath__39_I844 (.Y(N1814), .A0(N1737), .A1(N1734), .B0(N1736));
AOI21XL inst_blk01_cellmath__39_I848 (.Y(N1818), .A0(N1741), .A1(N1738), .B0(N1740));
NAND2XL inst_blk01_cellmath__39_I849 (.Y(N1819), .A(N1741), .B(N1739));
OAI21X2 inst_blk01_cellmath__39_I856 (.Y(N1826), .A0(N1819), .A1(N1814), .B0(N1818));
AOI21X2 inst_blk01_cellmath__39_I860 (.Y(N1830), .A0(N1745), .A1(N1742), .B0(N1744));
NAND2X1 inst_blk01_cellmath__39_I861 (.Y(N1831), .A(N1745), .B(N1743));
INVXL inst_blk01_cellmath__39_I1631 (.Y(N3055), .A(N1747));
AOI21X2 inst_blk01_cellmath__39_I864 (.Y(N1834), .A0(N1749), .A1(N1746), .B0(N1748));
NAND2X4 inst_blk01_cellmath__39_I865 (.Y(N1835), .A(N1749), .B(N1747));
OAI21X2 inst_blk01_cellmath__39_I872 (.Y(N1842), .A0(N1835), .A1(N1830), .B0(N1834));
NOR2X2 inst_blk01_cellmath__39_I873 (.Y(N1843), .A(N1835), .B(N1831));
AOI21X2 inst_blk01_cellmath__39_I876 (.Y(N1846), .A0(N1753), .A1(N1750), .B0(N1752));
NAND2X2 inst_blk01_cellmath__39_I877 (.Y(N1847), .A(N1753), .B(N1751));
INVXL inst_blk01_cellmath__39_I1641 (.Y(N3065), .A(N1755));
AOI21X4 inst_blk01_cellmath__39_I880 (.Y(N1850), .A0(N1757), .A1(N1754), .B0(N1756));
NAND2X4 inst_blk01_cellmath__39_I881 (.Y(N1851), .A(N1757), .B(N1755));
OAI21X4 inst_blk01_cellmath__39_I888 (.Y(N1858), .A0(N1851), .A1(N1846), .B0(N1850));
NOR2X4 inst_blk01_cellmath__39_I889 (.Y(N1859), .A(N1851), .B(N1847));
AOI21X4 inst_blk01_cellmath__39_I892 (.Y(N1862), .A0(N1761), .A1(N1758), .B0(N1760));
NAND2X4 inst_blk01_cellmath__39_I893 (.Y(N1863), .A(N1761), .B(N1759));
INVXL inst_blk01_cellmath__39_I1649 (.Y(N3073), .A(N1763));
AOI21X4 inst_blk01_cellmath__39_I896 (.Y(N1866), .A0(N1765), .A1(N1762), .B0(N1764));
NAND2X4 inst_blk01_cellmath__39_I897 (.Y(N1867), .A(N1765), .B(N1763));
OAI21X4 inst_blk01_cellmath__39_I904 (.Y(N1874), .A0(N1867), .A1(N1862), .B0(N1866));
NOR2X6 inst_blk01_cellmath__39_I905 (.Y(N1875), .A(N1867), .B(N1863));
AOI21X4 inst_blk01_cellmath__39_I908 (.Y(N1878), .A0(N1769), .A1(N1766), .B0(N1768));
NAND2X4 inst_blk01_cellmath__39_I909 (.Y(N1879), .A(N1769), .B(N1767));
INVXL inst_blk01_cellmath__39_I1659 (.Y(N3083), .A(N1771));
AOI21X4 inst_blk01_cellmath__39_I912 (.Y(N1882), .A0(N1773), .A1(N1770), .B0(N1772));
NAND2X6 inst_blk01_cellmath__39_I913 (.Y(N1883), .A(N1773), .B(N1771));
OAI21X4 inst_blk01_cellmath__39_I920 (.Y(N1890), .A0(N1883), .A1(N1878), .B0(N1882));
NOR2X6 inst_blk01_cellmath__39_I921 (.Y(N1891), .A(N1883), .B(N1879));
AOI21X4 inst_blk01_cellmath__39_I924 (.Y(N1894), .A0(N1777), .A1(N1774), .B0(N1776));
NAND2X4 inst_blk01_cellmath__39_I925 (.Y(N1895), .A(N1777), .B(N1775));
INVXL inst_blk01_cellmath__39_I1669 (.Y(N3093), .A(N1779));
AOI21X2 inst_blk01_cellmath__39_I928 (.Y(N1898), .A0(N1781), .A1(N1778), .B0(N1780));
NAND2X4 inst_blk01_cellmath__39_I929 (.Y(N1899), .A(N1781), .B(N1779));
OAI21X4 inst_blk01_cellmath__39_I936 (.Y(N1906), .A0(N1899), .A1(N1894), .B0(N1898));
NOR2X4 inst_blk01_cellmath__39_I937 (.Y(N1907), .A(N1899), .B(N1895));
AOI21X2 inst_blk01_cellmath__39_I940 (.Y(N1910), .A0(N1785), .A1(N1782), .B0(N1784));
NAND2X4 inst_blk01_cellmath__39_I941 (.Y(N1911), .A(N1785), .B(N1783));
INVXL inst_blk01_cellmath__39_I1677 (.Y(N3101), .A(N1787));
AOI21XL inst_blk01_cellmath__39_I944 (.Y(N1914), .A0(N1789), .A1(N1786), .B0(N1788));
NAND2X2 inst_blk01_cellmath__39_I945 (.Y(N1915), .A(N1789), .B(N1787));
OAI21X4 inst_blk01_cellmath__39_I952 (.Y(N1922), .A0(N1915), .A1(N1910), .B0(N1914));
NOR2X4 inst_blk01_cellmath__39_I953 (.Y(N1923), .A(N1915), .B(N1911));
AOI21X1 inst_blk01_cellmath__39_I956 (.Y(N1926), .A0(N1793), .A1(N1790), .B0(N1792));
NAND2X1 inst_blk01_cellmath__39_I957 (.Y(N1927), .A(N1793), .B(N1791));
INVXL inst_blk01_cellmath__39_I1685 (.Y(N3109), .A(N1795));
AOI21XL inst_blk01_cellmath__39_I960 (.Y(N1930), .A0(N1797), .A1(N1794), .B0(N1796));
NAND2XL inst_blk01_cellmath__39_I961 (.Y(N1931), .A(N1797), .B(N1795));
OAI21XL inst_blk01_cellmath__39_I968 (.Y(N1938), .A0(N1931), .A1(N1926), .B0(N1930));
NOR2XL inst_blk01_cellmath__39_I969 (.Y(N1939), .A(N1931), .B(N1927));
AOI21XL inst_blk01_cellmath__39_I972 (.Y(N1942), .A0(N1801), .A1(N1798), .B0(N1800));
NAND2XL inst_blk01_cellmath__39_I973 (.Y(N1943), .A(N1801), .B(N1799));
INVXL inst_blk01_cellmath__39_I1692 (.Y(N3116), .A(N1802));
INVXL inst_blk01_cellmath__39_I1693 (.Y(N3117), .A(N1803));
AOI21XL inst_blk01_cellmath__39_I976 (.Y(N1946), .A0(N1805), .A1(N1802), .B0(N1804));
NAND2XL inst_blk01_cellmath__39_I977 (.Y(N1947), .A(N1805), .B(N1803));
INVXL inst_blk01_cellmath__39_I1696 (.Y(N3120), .A(N1942));
INVXL inst_blk01_cellmath__39_I1697 (.Y(N3121), .A(N1943));
OAI21XL inst_blk01_cellmath__39_I982 (.Y(N1952), .A0(N3117), .A1(N1942), .B0(N3116));
NOR2XL inst_blk01_cellmath__39_I983 (.Y(N1953), .A(N3117), .B(N1943));
OAI21XL inst_blk01_cellmath__39_I984 (.Y(N1954), .A0(N1947), .A1(N1942), .B0(N1946));
NOR2XL inst_blk01_cellmath__39_I985 (.Y(N1955), .A(N1947), .B(N1943));
AOI21XL inst_blk01_cellmath__39_I994 (.Y(N1964), .A0(N1799), .A1(N1938), .B0(N1798));
AOI21XL inst_blk01_cellmath__39_I996 (.Y(N1966), .A0(N3121), .A1(N1938), .B0(N3120));
AOI21XL inst_blk01_cellmath__39_I998 (.Y(N1968), .A0(N1953), .A1(N1938), .B0(N1952));
AOI21XL inst_blk01_cellmath__39_I1004 (.Y(N1974), .A0(N1809), .A1(N1806), .B0(N1808));
NAND2XL inst_blk01_cellmath__39_I1005 (.Y(N1975), .A(N1809), .B(N1807));
INVXL inst_blk01_cellmath__39_I1709 (.Y(N3133), .A(N1811));
AO21XL inst_blk01_cellmath__39_I1823 (.Y(N3152), .A0(N1955), .A1(N1938), .B0(N1954));
AND2X1 inst_blk01_cellmath__39_I1824 (.Y(N3153), .A(N1939), .B(N1955));
INVXL inst_blk01_cellmath__39_I1730 (.Y(N3154), .A(N1826));
AOI21X2 inst_blk01_cellmath__39_I1032 (.Y(N2002), .A0(N1843), .A1(N1826), .B0(N1842));
AOI21X2 inst_blk01_cellmath__39_I1034 (.Y(N2004), .A0(N1859), .A1(N1842), .B0(N1858));
NAND2X2 inst_blk01_cellmath__39_I1035 (.Y(N2005), .A(N1859), .B(N1843));
AOI21X4 inst_blk01_cellmath__39_I1036 (.Y(N2006), .A0(N1875), .A1(N1858), .B0(N1874));
NAND2X4 inst_blk01_cellmath__39_I1037 (.Y(N2007), .A(N1875), .B(N1859));
AOI21X4 inst_blk01_cellmath__39_I1038 (.Y(N2008), .A0(N1891), .A1(N1874), .B0(N1890));
NAND2X4 inst_blk01_cellmath__39_I1039 (.Y(N2009), .A(N1891), .B(N1875));
AOI21X4 inst_blk01_cellmath__39_I1040 (.Y(N2010), .A0(N1907), .A1(N1890), .B0(N1906));
NAND2X4 inst_blk01_cellmath__39_I1041 (.Y(N2011), .A(N1907), .B(N1891));
AOI21X2 inst_blk01_cellmath__39_I1042 (.Y(N2012), .A0(N1923), .A1(N1906), .B0(N1922));
NAND2X2 inst_blk01_cellmath__39_I1043 (.Y(N2013), .A(N1923), .B(N1907));
AOI21X4 inst_blk01_cellmath__39_I1044 (.Y(N2014), .A0(N3153), .A1(N1922), .B0(N3152));
NAND2X4 inst_blk01_cellmath__39_I1045 (.Y(N2015), .A(N3153), .B(N1923));
INVXL inst_blk01_cellmath__39_I1731 (.Y(N3155), .A(N3154));
INVXL inst_blk01_cellmath__39_I1732 (.Y(N3156), .A(N2002));
OAI21X4 inst_blk01_cellmath__39_I1050 (.Y(N2020), .A0(N2005), .A1(N3154), .B0(N2004));
OAI21X4 inst_blk01_cellmath__39_I1052 (.Y(N2022), .A0(N2007), .A1(N2002), .B0(N2006));
OAI21X1 inst_blk01_cellmath__39_I1054 (.Y(N2024), .A0(N2009), .A1(N2004), .B0(N2008));
NOR2X1 inst_blk01_cellmath__39_I1055 (.Y(N2025), .A(N2009), .B(N2005));
OAI21X2 inst_blk01_cellmath__39_I1056 (.Y(N2026), .A0(N2011), .A1(N2006), .B0(N2010));
NOR2X1 inst_blk01_cellmath__39_I1057 (.Y(N2027), .A(N2011), .B(N2007));
OAI21X2 inst_blk01_cellmath__39_I1058 (.Y(N2028), .A0(N2013), .A1(N2008), .B0(N2012));
NOR2X2 inst_blk01_cellmath__39_I1059 (.Y(N2029), .A(N2013), .B(N2009));
OAI21X4 inst_blk01_cellmath__39_I1060 (.Y(N2030), .A0(N2015), .A1(N2010), .B0(N2014));
NOR2X2 inst_blk01_cellmath__39_I1061 (.Y(N2031), .A(N2015), .B(N2011));
INVXL inst_blk01_cellmath__39_I1733 (.Y(N3157), .A(N3155));
INVXL inst_blk01_cellmath__39_I1734 (.Y(N3158), .A(N3156));
INVXL inst_blk01_cellmath__39_I1735 (.Y(N3159), .A(N2020));
INVXL inst_blk01_cellmath__39_I1736 (.Y(N3160), .A(N2022));
AOI21X2 inst_blk01_cellmath__39_I1070 (.Y(N2040), .A0(N2025), .A1(N3155), .B0(N2024));
AOI21X2 inst_blk01_cellmath__39_I1072 (.Y(N2042), .A0(N2027), .A1(N3156), .B0(N2026));
AOI21X4 inst_blk01_cellmath__39_I1074 (.Y(N2044), .A0(N2029), .A1(N2020), .B0(N2028));
AOI21X4 inst_blk01_cellmath__39_I1076 (.Y(N2046), .A0(N2031), .A1(N2022), .B0(N2030));
NOR2BX1 andori2bb1_A_I3263 (.Y(N3245), .AN(N1739), .B(N1814));
NOR2XL andori2bb1_A_I1901 (.Y(N3165), .A(N3245), .B(N1738));
NOR2XL andori2bb1_A_I1902 (.Y(N3252), .A(N3055), .B(N1830));
NOR2XL andori2bb1_A_I1903 (.Y(N3170), .A(N3252), .B(N1746));
NOR2XL andori2bb1_A_I1904 (.Y(N3259), .A(N3065), .B(N1846));
NOR2XL andori2bb1_A_I1905 (.Y(N3176), .A(N3259), .B(N1754));
NOR2XL andori2bb1_A_I1908 (.Y(N3271), .A(N3073), .B(N1862));
NOR2XL andori2bb1_A_I1909 (.Y(N3182), .A(N3271), .B(N1762));
NOR2XL andori2bb1_A_I1910 (.Y(N3278), .A(N3083), .B(N1878));
NOR2XL andori2bb1_A_I1911 (.Y(N3188), .A(N3278), .B(N1770));
NOR2XL andori2bb1_A_I1912 (.Y(N3285), .A(N3093), .B(N1894));
NOR2XL andori2bb1_A_I1913 (.Y(N3194), .A(N3285), .B(N1778));
NOR2XL andori2bb1_A_I1914 (.Y(N3292), .A(N3101), .B(N1910));
NOR2XL andori2bb1_A_I1915 (.Y(N3200), .A(N3292), .B(N1786));
NOR2XL andori2bb1_A_I1916 (.Y(N3299), .A(N3109), .B(N1926));
NOR2XL andori2bb1_A_I1917 (.Y(N3206), .A(N3299), .B(N1794));
INVXL inst_blk01_cellmath__39_I1784 (.Y(N3208), .A(N1938));
NOR2XL andori2bb1_A_I1918 (.Y(N3306), .A(N3133), .B(N1974));
NOR2XL andori2bb1_A_I1919 (.Y(N3220), .A(N3306), .B(N1810));
OR2XL inst_blk01_cellmath__39_I1842 (.Y(N3221), .A(N3133), .B(N1975));
NAND2BXL inst_blk01_cellmath__39_I1184 (.Y(N2154), .AN(N1736), .B(N1737));
NAND2BXL inst_blk01_cellmath__39_I1187 (.Y(N2157), .AN(N1738), .B(N1739));
NAND2BXL inst_blk01_cellmath__39_I1190 (.Y(N2160), .AN(N1740), .B(N1741));
NAND2BXL inst_blk01_cellmath__39_I1193 (.Y(N2163), .AN(N1742), .B(N1743));
NAND2BXL inst_blk01_cellmath__39_I1196 (.Y(N2166), .AN(N1744), .B(N1745));
NAND2BXL inst_blk01_cellmath__39_I1199 (.Y(N2555), .AN(N1746), .B(N1747));
NAND2BXL inst_blk01_cellmath__39_I1202 (.Y(N2566), .AN(N1748), .B(N1749));
NAND2BXL inst_blk01_cellmath__39_I1205 (.Y(N2175), .AN(N1750), .B(N1751));
NAND2BXL inst_blk01_cellmath__39_I1208 (.Y(N2178), .AN(N1752), .B(N1753));
NAND2BXL inst_blk01_cellmath__39_I1211 (.Y(N2584), .AN(N1754), .B(N1755));
NAND2BXL inst_blk01_cellmath__39_I1214 (.Y(N2595), .AN(N1756), .B(N1757));
NAND2BXL inst_blk01_cellmath__39_I1217 (.Y(N2187), .AN(N1758), .B(N1759));
NAND2BXL inst_blk01_cellmath__39_I1220 (.Y(N2190), .AN(N1760), .B(N1761));
NAND2BXL inst_blk01_cellmath__39_I1223 (.Y(N2613), .AN(N1762), .B(N1763));
NAND2BXL inst_blk01_cellmath__39_I1226 (.Y(N2624), .AN(N1764), .B(N1765));
NAND2BXL inst_blk01_cellmath__39_I1229 (.Y(N2199), .AN(N1766), .B(N1767));
NAND2BXL inst_blk01_cellmath__39_I1232 (.Y(N2202), .AN(N1768), .B(N1769));
NAND2BXL inst_blk01_cellmath__39_I1235 (.Y(N2642), .AN(N1770), .B(N1771));
NAND2BXL inst_blk01_cellmath__39_I1238 (.Y(N2653), .AN(N1772), .B(N1773));
NAND2BXL inst_blk01_cellmath__39_I1241 (.Y(N2211), .AN(N1774), .B(N1775));
NAND2BXL inst_blk01_cellmath__39_I1244 (.Y(N2214), .AN(N1776), .B(N1777));
NAND2BXL inst_blk01_cellmath__39_I1247 (.Y(N2671), .AN(N1778), .B(N1779));
NAND2BXL inst_blk01_cellmath__39_I1250 (.Y(N2682), .AN(N1780), .B(N1781));
NAND2BXL inst_blk01_cellmath__39_I1253 (.Y(N2223), .AN(N1782), .B(N1783));
NAND2BXL inst_blk01_cellmath__39_I1256 (.Y(N2226), .AN(N1784), .B(N1785));
NAND2BXL inst_blk01_cellmath__39_I1259 (.Y(N2700), .AN(N1786), .B(N1787));
NAND2BXL inst_blk01_cellmath__39_I1262 (.Y(N2711), .AN(N1788), .B(N1789));
NAND2BXL inst_blk01_cellmath__39_I1265 (.Y(N2235), .AN(N1790), .B(N1791));
NAND2BXL inst_blk01_cellmath__39_I1268 (.Y(N2238), .AN(N1792), .B(N1793));
NAND2BXL inst_blk01_cellmath__39_I1271 (.Y(N2729), .AN(N1794), .B(N1795));
NAND2BXL inst_blk01_cellmath__39_I1274 (.Y(N2740), .AN(N1796), .B(N1797));
NAND2BXL inst_blk01_cellmath__39_I1277 (.Y(N2751), .AN(N1798), .B(N1799));
NAND2BXL inst_blk01_cellmath__39_I1280 (.Y(N2762), .AN(N1800), .B(N1801));
NAND2BXL inst_blk01_cellmath__39_I1283 (.Y(N2773), .AN(N1802), .B(N1803));
NAND2BXL inst_blk01_cellmath__39_I1286 (.Y(N2784), .AN(N1804), .B(N1805));
NAND2BXL inst_blk01_cellmath__39_I1289 (.Y(N2259), .AN(N1806), .B(N1807));
NAND2BXL inst_blk01_cellmath__39_I1292 (.Y(N2262), .AN(N1808), .B(N1809));
NAND2BXL inst_blk01_cellmath__39_I1295 (.Y(N2802), .AN(N1810), .B(N1811));
XOR2XL inst_blk01_cellmath__39_I1843 (.Y(inst_blk01_cellmath__39_out0[16]), .A(N1734), .B(N2154));
XNOR2X1 inst_blk01_cellmath__39_I1298 (.Y(inst_blk01_cellmath__39_out0[17]), .A(N1814), .B(N2157));
XNOR2X1 inst_blk01_cellmath__39_I1299 (.Y(inst_blk01_cellmath__39_out0[18]), .A(N3165), .B(N2160));
XNOR2X1 inst_blk01_cellmath__39_I1300 (.Y(inst_blk01_cellmath__39_out0[19]), .A(N3157), .B(N2163));
XNOR2X1 inst_blk01_cellmath__39_I1301 (.Y(inst_blk01_cellmath__39_out0[23]), .A(N3158), .B(N2175));
XNOR2X1 inst_blk01_cellmath__39_I1302 (.Y(inst_blk01_cellmath__39_out0[27]), .A(N3159), .B(N2187));
XNOR2X1 inst_blk01_cellmath__39_I1303 (.Y(inst_blk01_cellmath__39_out0[31]), .A(N3160), .B(N2199));
XNOR2XL inst_blk01_cellmath__39_I1304 (.Y(inst_blk01_cellmath__39_out0[35]), .A(N2040), .B(N2211));
XNOR2XL inst_blk01_cellmath__39_I1305 (.Y(inst_blk01_cellmath__39_out0[39]), .A(N2042), .B(N2223));
XNOR2XL inst_blk01_cellmath__39_I1306 (.Y(inst_blk01_cellmath__39_out0[43]), .A(N2044), .B(N2235));
XNOR2X1 inst_blk01_cellmath__39_I1307 (.Y(inst_blk01_cellmath__39_out0[51]), .A(N2046), .B(N2259));
XOR2XL node_cs_reduced_ii_local_A_I1844 (.Y(N2279), .A(N2166), .B(N1743));
XOR2XL node_cs_reduced_ii_local_A_I1845 (.Y(N2278), .A(N2166), .B(N1742));
MX2XL inst_blk01_cellmath__39_I1309 (.Y(inst_blk01_cellmath__39_out0[20]), .A(N2279), .B(N2278), .S0(N3157));
XOR2XL node_cs_ii_local_alt_A_I1429 (.Y(N2281), .A(N2555), .B(N1830));
NAND2XL node_cs_ii_local_alt_A_I1430 (.Y(N2553), .A(N1831), .B(N1830));
XNOR2X1 node_cs_ii_local_alt_A_I1431 (.Y(N2282), .A(N2555), .B(N2553));
MXI2XL inst_blk01_cellmath__39_I1311 (.Y(inst_blk01_cellmath__39_out0[21]), .A(N2282), .B(N2281), .S0(N3157));
XOR2XL node_cs_ii_local_alt_A_I1433 (.Y(N2284), .A(N2566), .B(N3170));
OAI21XL node_cs_ii_local_alt_A_I1846 (.Y(N2564), .A0(N3055), .A1(N1831), .B0(N3170));
XNOR2X1 node_cs_ii_local_alt_A_I1435 (.Y(N2285), .A(N2566), .B(N2564));
MXI2XL inst_blk01_cellmath__39_I1313 (.Y(inst_blk01_cellmath__39_out0[22]), .A(N2285), .B(N2284), .S0(N3157));
XOR2XL node_cs_reduced_ii_local_A_I1847 (.Y(N2288), .A(N2178), .B(N1751));
XOR2XL node_cs_reduced_ii_local_A_I1848 (.Y(N2287), .A(N2178), .B(N1750));
MX2XL inst_blk01_cellmath__39_I1315 (.Y(inst_blk01_cellmath__39_out0[24]), .A(N2288), .B(N2287), .S0(N3158));
XOR2XL node_cs_ii_local_alt_A_I1439 (.Y(N2290), .A(N2584), .B(N1846));
NAND2XL node_cs_ii_local_alt_A_I1440 (.Y(N2582), .A(N1847), .B(N1846));
XNOR2X1 node_cs_ii_local_alt_A_I1441 (.Y(N2291), .A(N2584), .B(N2582));
MXI2XL inst_blk01_cellmath__39_I1317 (.Y(inst_blk01_cellmath__39_out0[25]), .A(N2291), .B(N2290), .S0(N3158));
XOR2XL node_cs_ii_local_alt_A_I1443 (.Y(N2293), .A(N2595), .B(N3176));
OAI21XL node_cs_ii_local_alt_A_I1849 (.Y(N2593), .A0(N3065), .A1(N1847), .B0(N3176));
XNOR2X1 node_cs_ii_local_alt_A_I1445 (.Y(N2294), .A(N2595), .B(N2593));
MXI2XL inst_blk01_cellmath__39_I1319 (.Y(inst_blk01_cellmath__39_out0[26]), .A(N2294), .B(N2293), .S0(N3158));
XOR2XL node_cs_reduced_ii_local_A_I1850 (.Y(N2297), .A(N2190), .B(N1759));
XOR2XL node_cs_reduced_ii_local_A_I1851 (.Y(N2296), .A(N2190), .B(N1758));
MX2XL inst_blk01_cellmath__39_I1321 (.Y(inst_blk01_cellmath__39_out0[28]), .A(N2297), .B(N2296), .S0(N3159));
XOR2XL node_cs_ii_local_alt_A_I1449 (.Y(N2299), .A(N2613), .B(N1862));
NAND2XL node_cs_ii_local_alt_A_I1450 (.Y(N2611), .A(N1863), .B(N1862));
XNOR2X1 node_cs_ii_local_alt_A_I1451 (.Y(N2300), .A(N2613), .B(N2611));
MXI2XL inst_blk01_cellmath__39_I1323 (.Y(inst_blk01_cellmath__39_out0[29]), .A(N2300), .B(N2299), .S0(N3159));
XOR2XL node_cs_ii_local_alt_A_I1453 (.Y(N2302), .A(N2624), .B(N3182));
OAI21XL node_cs_ii_local_alt_A_I1852 (.Y(N2622), .A0(N3073), .A1(N1863), .B0(N3182));
XNOR2X1 node_cs_ii_local_alt_A_I1455 (.Y(N2303), .A(N2624), .B(N2622));
MXI2XL inst_blk01_cellmath__39_I1325 (.Y(inst_blk01_cellmath__39_out0[30]), .A(N2303), .B(N2302), .S0(N3159));
XOR2XL node_cs_reduced_ii_local_A_I1853 (.Y(N2306), .A(N2202), .B(N1767));
XOR2XL node_cs_reduced_ii_local_A_I1854 (.Y(N2305), .A(N2202), .B(N1766));
MX2XL inst_blk01_cellmath__39_I1327 (.Y(inst_blk01_cellmath__39_out0[32]), .A(N2306), .B(N2305), .S0(N3160));
XOR2XL node_cs_ii_local_alt_A_I1459 (.Y(N2308), .A(N2642), .B(N1878));
NAND2XL node_cs_ii_local_alt_A_I1460 (.Y(N2640), .A(N1879), .B(N1878));
XNOR2X1 node_cs_ii_local_alt_A_I1461 (.Y(N2309), .A(N2642), .B(N2640));
MXI2XL inst_blk01_cellmath__39_I1329 (.Y(inst_blk01_cellmath__39_out0[33]), .A(N2309), .B(N2308), .S0(N3160));
XOR2XL node_cs_ii_local_alt_A_I1463 (.Y(N2311), .A(N2653), .B(N3188));
OAI21XL node_cs_ii_local_alt_A_I1887 (.Y(N2651), .A0(N3083), .A1(N1879), .B0(N3188));
XNOR2X1 node_cs_ii_local_alt_A_I1465 (.Y(N2312), .A(N2653), .B(N2651));
MXI2XL inst_blk01_cellmath__39_I1331 (.Y(inst_blk01_cellmath__39_out0[34]), .A(N2312), .B(N2311), .S0(N3160));
XOR2XL node_cs_reduced_ii_local_A_I1856 (.Y(N2315), .A(N2214), .B(N1775));
XOR2XL node_cs_reduced_ii_local_A_I1857 (.Y(N2314), .A(N2214), .B(N1774));
MX2XL inst_blk01_cellmath__39_I1333 (.Y(inst_blk01_cellmath__39_out0[36]), .A(N2315), .B(N2314), .S0(N2040));
XOR2XL node_cs_ii_local_alt_A_I1469 (.Y(N2317), .A(N2671), .B(N1894));
NAND2XL node_cs_ii_local_alt_A_I1470 (.Y(N2669), .A(N1895), .B(N1894));
XNOR2X1 node_cs_ii_local_alt_A_I1471 (.Y(N2318), .A(N2671), .B(N2669));
MXI2XL inst_blk01_cellmath__39_I1335 (.Y(inst_blk01_cellmath__39_out0[37]), .A(N2318), .B(N2317), .S0(N2040));
XOR2XL node_cs_ii_local_alt_A_I1473 (.Y(N2320), .A(N2682), .B(N3194));
OAI21XL node_cs_ii_local_alt_A_I1858 (.Y(N2680), .A0(N3093), .A1(N1895), .B0(N3194));
XNOR2X1 node_cs_ii_local_alt_A_I1475 (.Y(N2321), .A(N2682), .B(N2680));
MXI2XL inst_blk01_cellmath__39_I1337 (.Y(inst_blk01_cellmath__39_out0[38]), .A(N2321), .B(N2320), .S0(N2040));
XOR2XL node_cs_reduced_ii_local_A_I1859 (.Y(N2324), .A(N2226), .B(N1783));
XOR2XL node_cs_reduced_ii_local_A_I1860 (.Y(N2323), .A(N2226), .B(N1782));
MX2XL inst_blk01_cellmath__39_I1339 (.Y(inst_blk01_cellmath__39_out0[40]), .A(N2324), .B(N2323), .S0(N2042));
XOR2XL node_cs_ii_local_alt_A_I1479 (.Y(N2326), .A(N2700), .B(N1910));
NAND2XL node_cs_ii_local_alt_A_I1480 (.Y(N2698), .A(N1911), .B(N1910));
XNOR2X1 node_cs_ii_local_alt_A_I1481 (.Y(N2327), .A(N2700), .B(N2698));
MXI2XL inst_blk01_cellmath__39_I1341 (.Y(inst_blk01_cellmath__39_out0[41]), .A(N2327), .B(N2326), .S0(N2042));
XOR2XL node_cs_ii_local_alt_A_I1483 (.Y(N2329), .A(N2711), .B(N3200));
OAI21XL node_cs_ii_local_alt_A_I1861 (.Y(N2709), .A0(N3101), .A1(N1911), .B0(N3200));
XNOR2X1 node_cs_ii_local_alt_A_I1485 (.Y(N2330), .A(N2711), .B(N2709));
MXI2XL inst_blk01_cellmath__39_I1343 (.Y(inst_blk01_cellmath__39_out0[42]), .A(N2330), .B(N2329), .S0(N2042));
XOR2XL node_cs_reduced_ii_local_A_I1862 (.Y(N2333), .A(N2238), .B(N1791));
XOR2XL node_cs_reduced_ii_local_A_I1863 (.Y(N2332), .A(N2238), .B(N1790));
MX2XL inst_blk01_cellmath__39_I1345 (.Y(inst_blk01_cellmath__39_out0[44]), .A(N2333), .B(N2332), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1489 (.Y(N2335), .A(N2729), .B(N1926));
NAND2XL node_cs_ii_local_alt_A_I1490 (.Y(N2727), .A(N1927), .B(N1926));
XNOR2X1 node_cs_ii_local_alt_A_I1491 (.Y(N2336), .A(N2729), .B(N2727));
MXI2XL inst_blk01_cellmath__39_I1347 (.Y(inst_blk01_cellmath__39_out0[45]), .A(N2336), .B(N2335), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1493 (.Y(N2338), .A(N2740), .B(N3206));
OAI21XL node_cs_ii_local_alt_A_I1864 (.Y(N2738), .A0(N3109), .A1(N1927), .B0(N3206));
XNOR2X1 node_cs_ii_local_alt_A_I1495 (.Y(N2339), .A(N2740), .B(N2738));
MXI2XL inst_blk01_cellmath__39_I1349 (.Y(inst_blk01_cellmath__39_out0[46]), .A(N2339), .B(N2338), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1497 (.Y(N2341), .A(N2751), .B(N3208));
NAND2BXL node_cs_ii_local_alt_A_I1865 (.Y(N2749), .AN(N1939), .B(N3208));
XNOR2X1 node_cs_ii_local_alt_A_I1499 (.Y(N2342), .A(N2751), .B(N2749));
MXI2XL inst_blk01_cellmath__39_I1351 (.Y(inst_blk01_cellmath__39_out0[47]), .A(N2342), .B(N2341), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1501 (.Y(N2344), .A(N2762), .B(N1964));
OAI2BB1X1 node_cs_ii_local_alt_A_I1866 (.Y(N2760), .A0N(N1799), .A1N(N1939), .B0(N1964));
XNOR2X1 node_cs_ii_local_alt_A_I1503 (.Y(N2345), .A(N2762), .B(N2760));
MXI2XL inst_blk01_cellmath__39_I1353 (.Y(inst_blk01_cellmath__39_out0[48]), .A(N2345), .B(N2344), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1505 (.Y(N2347), .A(N2773), .B(N1966));
OAI2BB1X1 node_cs_ii_local_alt_A_I1867 (.Y(N2771), .A0N(N3121), .A1N(N1939), .B0(N1966));
XNOR2X1 node_cs_ii_local_alt_A_I1507 (.Y(N2348), .A(N2773), .B(N2771));
MXI2XL inst_blk01_cellmath__39_I1355 (.Y(inst_blk01_cellmath__39_out0[49]), .A(N2348), .B(N2347), .S0(N2044));
XOR2XL node_cs_ii_local_alt_A_I1509 (.Y(N2350), .A(N2784), .B(N1968));
OAI2BB1X1 node_cs_ii_local_alt_A_I1868 (.Y(N2782), .A0N(N1953), .A1N(N1939), .B0(N1968));
XNOR2X1 node_cs_ii_local_alt_A_I1511 (.Y(N2351), .A(N2784), .B(N2782));
MXI2XL inst_blk01_cellmath__39_I1357 (.Y(inst_blk01_cellmath__39_out0[50]), .A(N2351), .B(N2350), .S0(N2044));
XOR2XL node_cs_reduced_ii_local_A_I1869 (.Y(N2354), .A(N2262), .B(N1807));
XOR2XL node_cs_reduced_ii_local_A_I1870 (.Y(N2353), .A(N2262), .B(N1806));
MX2XL inst_blk01_cellmath__39_I1359 (.Y(inst_blk01_cellmath__39_out0[52]), .A(N2354), .B(N2353), .S0(N2046));
XOR2XL node_cs_ii_local_alt_A_I1515 (.Y(N2356), .A(N2802), .B(N1974));
NAND2XL node_cs_ii_local_alt_A_I1516 (.Y(N2800), .A(N1975), .B(N1974));
XNOR2X1 node_cs_ii_local_alt_A_I1517 (.Y(N2357), .A(N2802), .B(N2800));
MXI2XL inst_blk01_cellmath__39_I1361 (.Y(inst_blk01_cellmath__39_out0[53]), .A(N2357), .B(N2356), .S0(N2046));
OA21X1 inst_blk01_cellmath__39_I1540 (.Y(inst_blk01_cellmath__39_out0[55]), .A0(N3221), .A1(N2046), .B0(N3220));
INVXL inst_blk01_cellmath__39_I1798 (.Y(inst_blk01_cellmath__39_out0[54]), .A(inst_blk01_cellmath__39_out0[55]));
assign inst_blk01_cellmath__39_out0[0] = 1'B0;
endmodule

module cynw_cm_float_sin_inst_cellmath__42_0_bdw1946085813_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0
	); /* architecture "gate_level" */ 
output [5:0] inst_cellmath__42_0_out0;
input [5:0] inst_cellmath__42_0_in0;
wire N25,N27,N49,N150,N160,N167;
INVX1 inst_cellmath__42_0_I5 (.Y(inst_cellmath__42_0_out0[0]), .A(inst_cellmath__42_0_in0[0]));
INVXL inst_cellmath__42_0_I80 (.Y(N150), .A(inst_cellmath__42_0_in0[1]));
INVXL inst_cellmath__42_0_I7 (.Y(N25), .A(inst_cellmath__42_0_in0[2]));
INVXL inst_cellmath__42_0_I8 (.Y(N27), .A(inst_cellmath__42_0_in0[3]));
OAI21XL inst_cellmath__42_0_I24 (.Y(N49), .A0(N25), .A1(N150), .B0(N27));
INVXL inst_cellmath__42_0_I86 (.Y(inst_cellmath__42_0_out0[1]), .A(N150));
MXI2XL inst_cellmath__42_0_I67 (.Y(inst_cellmath__42_0_out0[2]), .A(N150), .B(inst_cellmath__42_0_out0[1]), .S0(N25));
NOR2XL node_cs_const1_cs_A_I94 (.Y(N160), .A(N25), .B(N150));
XNOR2X1 node_cs_const1_cs_A_I95 (.Y(inst_cellmath__42_0_out0[3]), .A(N27), .B(N160));
XOR2XL inst_cellmath__42_0_I91 (.Y(inst_cellmath__42_0_out0[4]), .A(N49), .B(inst_cellmath__42_0_in0[4]));
NOR2XL node_cs_const1_cs_A_I96 (.Y(N167), .A(inst_cellmath__42_0_in0[4]), .B(N49));
XNOR2X1 node_cs_const1_cs_A_I97 (.Y(inst_cellmath__42_0_out0[5]), .A(inst_cellmath__42_0_in0[5]), .B(N167));
endmodule

module cynw_cm_float_sin_inst_cellmath__48_bdw1946085813_bdw (
	inst_cellmath__48_out0,
	inst_cellmath__48_in0,
	inst_cellmath__48_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__48_out0;
input [5:0] inst_cellmath__48_in0;
input [55:26] inst_cellmath__48_in1;
wire N65,N66,N67,N68,N69,N70,N71 
	,N72,N73,N74,N75,N76,N77,N78,N79 
	,N80,N81,N82,N83,N84,N85,N86,N87 
	,N88,N89,N90,N91,N92,N93,N94,N130 
	,N131,N132,N133,N134,N135,N136,N137,N138 
	,N139,N140,N141,N142,N143,N144,N145,N146 
	,N147,N148,N149,N150,N151,N152,N153,N154 
	,N155,N156,N157,N158,N160,N196,N197,N198 
	,N199,N200,N201,N202,N203,N204,N205,N206 
	,N207,N208,N209,N210,N211,N212,N213,N214 
	,N215,N216,N217,N218,N219,N220,N221,N222 
	,N224,N226,N228,N264,N265,N266,N267,N268 
	,N269,N270,N271,N272,N273,N274,N275,N276 
	,N277,N278,N280,N282,N284,N286,N288,N290 
	,N292,N294,N296,N298,N300,N302,N304,N306 
	,N308,N344,N345,N346,N347,N348,N349,N350 
	,N351,N352,N353,N354,N355,N356,N357,N358 
	,N359,N360,N361,N362,N363,N364,N365,N366 
	,N368,N370,N508,N509,N510,N511,N512,N513 
	,N514,N515,N516,N517,N518,N519,N520,N521 
	,N522,N523,N524,N525,N526,N527,N528,N529 
	,N530,N531,N532,N533,N534,N535,N536,N537 
	,N538,N539,N540,N541,N542,N543,N544,N545 
	,N546,N547,N548,N549,N550,N551,N552,N553 
	,N554,N555;
INVXL inst_cellmath__48_I384 (.Y(N508), .A(inst_cellmath__48_in0[0]));
INVXL inst_cellmath__48_I385 (.Y(N509), .A(N508));
INVXL inst_cellmath__48_I391 (.Y(N515), .A(N509));
INVXL inst_cellmath__48_I390 (.Y(N514), .A(N509));
INVXL inst_cellmath__48_I389 (.Y(N513), .A(N509));
INVXL inst_cellmath__48_I388 (.Y(N512), .A(N509));
INVXL inst_cellmath__48_I387 (.Y(N511), .A(N509));
INVXL inst_cellmath__48_I386 (.Y(N510), .A(N509));
MXI2XL inst_cellmath__48_I2 (.Y(N65), .A(inst_cellmath__48_in1[27]), .B(inst_cellmath__48_in1[26]), .S0(N515));
MXI2XL inst_cellmath__48_I3 (.Y(N66), .A(inst_cellmath__48_in1[28]), .B(inst_cellmath__48_in1[27]), .S0(N515));
MXI2XL inst_cellmath__48_I4 (.Y(N67), .A(inst_cellmath__48_in1[29]), .B(inst_cellmath__48_in1[28]), .S0(N515));
MXI2XL inst_cellmath__48_I5 (.Y(N68), .A(inst_cellmath__48_in1[30]), .B(inst_cellmath__48_in1[29]), .S0(N515));
MXI2XL inst_cellmath__48_I6 (.Y(N69), .A(inst_cellmath__48_in1[31]), .B(inst_cellmath__48_in1[30]), .S0(N515));
MXI2XL inst_cellmath__48_I7 (.Y(N70), .A(inst_cellmath__48_in1[32]), .B(inst_cellmath__48_in1[31]), .S0(N514));
MXI2XL inst_cellmath__48_I8 (.Y(N71), .A(inst_cellmath__48_in1[33]), .B(inst_cellmath__48_in1[32]), .S0(N514));
MXI2XL inst_cellmath__48_I9 (.Y(N72), .A(inst_cellmath__48_in1[34]), .B(inst_cellmath__48_in1[33]), .S0(N514));
MXI2XL inst_cellmath__48_I10 (.Y(N73), .A(inst_cellmath__48_in1[35]), .B(inst_cellmath__48_in1[34]), .S0(N514));
MXI2XL inst_cellmath__48_I11 (.Y(N74), .A(inst_cellmath__48_in1[36]), .B(inst_cellmath__48_in1[35]), .S0(N514));
MXI2XL inst_cellmath__48_I12 (.Y(N75), .A(inst_cellmath__48_in1[37]), .B(inst_cellmath__48_in1[36]), .S0(N513));
MXI2XL inst_cellmath__48_I13 (.Y(N76), .A(inst_cellmath__48_in1[38]), .B(inst_cellmath__48_in1[37]), .S0(N513));
MXI2XL inst_cellmath__48_I14 (.Y(N77), .A(inst_cellmath__48_in1[39]), .B(inst_cellmath__48_in1[38]), .S0(N513));
MXI2XL inst_cellmath__48_I15 (.Y(N78), .A(inst_cellmath__48_in1[40]), .B(inst_cellmath__48_in1[39]), .S0(N513));
MXI2XL inst_cellmath__48_I16 (.Y(N79), .A(inst_cellmath__48_in1[41]), .B(inst_cellmath__48_in1[40]), .S0(N513));
MXI2XL inst_cellmath__48_I17 (.Y(N80), .A(inst_cellmath__48_in1[42]), .B(inst_cellmath__48_in1[41]), .S0(N512));
MXI2XL inst_cellmath__48_I18 (.Y(N81), .A(inst_cellmath__48_in1[43]), .B(inst_cellmath__48_in1[42]), .S0(N512));
MXI2XL inst_cellmath__48_I19 (.Y(N82), .A(inst_cellmath__48_in1[44]), .B(inst_cellmath__48_in1[43]), .S0(N512));
MXI2XL inst_cellmath__48_I20 (.Y(N83), .A(inst_cellmath__48_in1[45]), .B(inst_cellmath__48_in1[44]), .S0(N512));
MXI2XL inst_cellmath__48_I21 (.Y(N84), .A(inst_cellmath__48_in1[46]), .B(inst_cellmath__48_in1[45]), .S0(N512));
MXI2XL inst_cellmath__48_I22 (.Y(N85), .A(inst_cellmath__48_in1[47]), .B(inst_cellmath__48_in1[46]), .S0(N511));
MXI2XL inst_cellmath__48_I23 (.Y(N86), .A(inst_cellmath__48_in1[48]), .B(inst_cellmath__48_in1[47]), .S0(N511));
MXI2X1 inst_cellmath__48_I24 (.Y(N87), .A(inst_cellmath__48_in1[49]), .B(inst_cellmath__48_in1[48]), .S0(N511));
MXI2X1 inst_cellmath__48_I25 (.Y(N88), .A(inst_cellmath__48_in1[50]), .B(inst_cellmath__48_in1[49]), .S0(N511));
MXI2XL inst_cellmath__48_I26 (.Y(N89), .A(inst_cellmath__48_in1[51]), .B(inst_cellmath__48_in1[50]), .S0(N511));
MXI2XL inst_cellmath__48_I27 (.Y(N90), .A(inst_cellmath__48_in1[52]), .B(inst_cellmath__48_in1[51]), .S0(N510));
MXI2XL inst_cellmath__48_I28 (.Y(N91), .A(inst_cellmath__48_in1[53]), .B(inst_cellmath__48_in1[52]), .S0(N510));
MXI2XL inst_cellmath__48_I29 (.Y(N92), .A(inst_cellmath__48_in1[54]), .B(inst_cellmath__48_in1[53]), .S0(N510));
MXI2XL inst_cellmath__48_I30 (.Y(N93), .A(inst_cellmath__48_in1[55]), .B(inst_cellmath__48_in1[54]), .S0(N510));
NAND2XL inst_cellmath__48_I31 (.Y(N94), .A(inst_cellmath__48_in1[55]), .B(N510));
INVXL inst_cellmath__48_I392 (.Y(N516), .A(inst_cellmath__48_in0[1]));
INVXL inst_cellmath__48_I398 (.Y(N522), .A(N516));
INVXL inst_cellmath__48_I397 (.Y(N521), .A(N516));
INVXL inst_cellmath__48_I396 (.Y(N520), .A(N516));
INVXL inst_cellmath__48_I395 (.Y(N519), .A(N516));
INVXL inst_cellmath__48_I394 (.Y(N518), .A(N516));
INVXL inst_cellmath__48_I393 (.Y(N517), .A(N516));
MXI2XL inst_cellmath__48_I66 (.Y(N130), .A(N65), .B(N67), .S0(N522));
MXI2XL inst_cellmath__48_I67 (.Y(N131), .A(N66), .B(N68), .S0(N522));
MXI2XL inst_cellmath__48_I68 (.Y(N132), .A(N67), .B(N69), .S0(N522));
MXI2XL inst_cellmath__48_I69 (.Y(N133), .A(N68), .B(N70), .S0(N522));
MXI2XL inst_cellmath__48_I70 (.Y(N134), .A(N69), .B(N71), .S0(N522));
MXI2XL inst_cellmath__48_I71 (.Y(N135), .A(N70), .B(N72), .S0(N521));
MXI2XL inst_cellmath__48_I72 (.Y(N136), .A(N71), .B(N73), .S0(N521));
MXI2XL inst_cellmath__48_I73 (.Y(N137), .A(N72), .B(N74), .S0(N521));
MXI2XL inst_cellmath__48_I74 (.Y(N138), .A(N73), .B(N75), .S0(N521));
MXI2XL inst_cellmath__48_I75 (.Y(N139), .A(N74), .B(N76), .S0(N521));
MXI2XL inst_cellmath__48_I76 (.Y(N140), .A(N75), .B(N77), .S0(N520));
MXI2XL inst_cellmath__48_I77 (.Y(N141), .A(N76), .B(N78), .S0(N520));
MXI2XL inst_cellmath__48_I78 (.Y(N142), .A(N77), .B(N79), .S0(N520));
MXI2XL inst_cellmath__48_I79 (.Y(N143), .A(N78), .B(N80), .S0(N520));
MXI2XL inst_cellmath__48_I80 (.Y(N144), .A(N79), .B(N81), .S0(N520));
MXI2XL inst_cellmath__48_I81 (.Y(N145), .A(N80), .B(N82), .S0(N519));
MXI2XL inst_cellmath__48_I82 (.Y(N146), .A(N81), .B(N83), .S0(N519));
MXI2XL inst_cellmath__48_I83 (.Y(N147), .A(N82), .B(N84), .S0(N519));
MXI2XL inst_cellmath__48_I84 (.Y(N148), .A(N83), .B(N85), .S0(N519));
MXI2XL inst_cellmath__48_I85 (.Y(N149), .A(N84), .B(N86), .S0(N519));
MXI2X1 inst_cellmath__48_I86 (.Y(N150), .A(N85), .B(N87), .S0(N518));
MXI2XL inst_cellmath__48_I87 (.Y(N151), .A(N86), .B(N88), .S0(N518));
MXI2X1 inst_cellmath__48_I88 (.Y(N152), .A(N87), .B(N89), .S0(N518));
MXI2X1 inst_cellmath__48_I89 (.Y(N153), .A(N88), .B(N90), .S0(N518));
MXI2X1 inst_cellmath__48_I90 (.Y(N154), .A(N89), .B(N91), .S0(N518));
MXI2XL inst_cellmath__48_I91 (.Y(N155), .A(N90), .B(N92), .S0(N517));
MXI2XL inst_cellmath__48_I92 (.Y(N156), .A(N91), .B(N93), .S0(N517));
MXI2X1 inst_cellmath__48_I93 (.Y(N157), .A(N92), .B(N94), .S0(N517));
NOR2XL inst_cellmath__48_I94 (.Y(N158), .A(N93), .B(N517));
NOR2XL inst_cellmath__48_I95 (.Y(N160), .A(N94), .B(N517));
INVXL inst_cellmath__48_I399 (.Y(N523), .A(inst_cellmath__48_in0[2]));
INVXL inst_cellmath__48_I400 (.Y(N524), .A(N523));
INVXL inst_cellmath__48_I406 (.Y(N530), .A(N524));
INVXL inst_cellmath__48_I405 (.Y(N529), .A(N524));
INVXL inst_cellmath__48_I404 (.Y(N528), .A(N524));
INVXL inst_cellmath__48_I403 (.Y(N527), .A(N524));
INVXL inst_cellmath__48_I402 (.Y(N526), .A(N524));
INVXL inst_cellmath__48_I401 (.Y(N525), .A(N524));
MXI2XL inst_cellmath__48_I130 (.Y(N196), .A(N134), .B(N130), .S0(N530));
MXI2XL inst_cellmath__48_I131 (.Y(N197), .A(N135), .B(N131), .S0(N530));
MXI2XL inst_cellmath__48_I132 (.Y(N198), .A(N136), .B(N132), .S0(N530));
MXI2XL inst_cellmath__48_I133 (.Y(N199), .A(N137), .B(N133), .S0(N530));
MXI2XL inst_cellmath__48_I134 (.Y(N200), .A(N138), .B(N134), .S0(N530));
MXI2XL inst_cellmath__48_I135 (.Y(N201), .A(N139), .B(N135), .S0(N529));
MXI2XL inst_cellmath__48_I136 (.Y(N202), .A(N140), .B(N136), .S0(N529));
MXI2XL inst_cellmath__48_I137 (.Y(N203), .A(N141), .B(N137), .S0(N529));
MXI2XL inst_cellmath__48_I138 (.Y(N204), .A(N142), .B(N138), .S0(N529));
MXI2XL inst_cellmath__48_I139 (.Y(N205), .A(N143), .B(N139), .S0(N529));
MXI2XL inst_cellmath__48_I140 (.Y(N206), .A(N144), .B(N140), .S0(N528));
MXI2XL inst_cellmath__48_I141 (.Y(N207), .A(N145), .B(N141), .S0(N528));
MXI2XL inst_cellmath__48_I142 (.Y(N208), .A(N146), .B(N142), .S0(N528));
MXI2XL inst_cellmath__48_I143 (.Y(N209), .A(N147), .B(N143), .S0(N528));
MXI2XL inst_cellmath__48_I144 (.Y(N210), .A(N148), .B(N144), .S0(N528));
MXI2XL inst_cellmath__48_I145 (.Y(N211), .A(N149), .B(N145), .S0(N527));
MXI2XL inst_cellmath__48_I146 (.Y(N212), .A(N150), .B(N146), .S0(N527));
MXI2X1 inst_cellmath__48_I147 (.Y(N213), .A(N151), .B(N147), .S0(N527));
MXI2X1 inst_cellmath__48_I148 (.Y(N214), .A(N152), .B(N148), .S0(N527));
MXI2XL inst_cellmath__48_I149 (.Y(N215), .A(N153), .B(N149), .S0(N527));
MXI2XL inst_cellmath__48_I150 (.Y(N216), .A(N154), .B(N150), .S0(N526));
MXI2XL inst_cellmath__48_I151 (.Y(N217), .A(N155), .B(N151), .S0(N526));
MXI2X1 inst_cellmath__48_I152 (.Y(N218), .A(N156), .B(N152), .S0(N526));
MXI2X1 inst_cellmath__48_I153 (.Y(N219), .A(N157), .B(N153), .S0(N526));
MXI2X1 inst_cellmath__48_I154 (.Y(N220), .A(N158), .B(N154), .S0(N526));
MXI2X1 inst_cellmath__48_I155 (.Y(N221), .A(N160), .B(N155), .S0(N525));
NAND2XL inst_cellmath__48_I156 (.Y(N222), .A(N156), .B(N525));
NAND2XL inst_cellmath__48_I157 (.Y(N224), .A(N157), .B(N525));
NAND2XL inst_cellmath__48_I158 (.Y(N226), .A(N158), .B(N525));
NAND2XL inst_cellmath__48_I159 (.Y(N228), .A(N160), .B(N525));
INVXL inst_cellmath__48_I407 (.Y(N531), .A(inst_cellmath__48_in0[4]));
INVXL inst_cellmath__48_I408 (.Y(N532), .A(N531));
INVXL inst_cellmath__48_I415 (.Y(N539), .A(N532));
INVXL inst_cellmath__48_I409 (.Y(N533), .A(N532));
INVXL inst_cellmath__48_I416 (.Y(N540), .A(N539));
INVXL inst_cellmath__48_I414 (.Y(N538), .A(N533));
INVXL inst_cellmath__48_I413 (.Y(N537), .A(N533));
INVXL inst_cellmath__48_I412 (.Y(N536), .A(N533));
INVXL inst_cellmath__48_I411 (.Y(N535), .A(N533));
INVXL inst_cellmath__48_I410 (.Y(N534), .A(N533));
MXI2XL inst_cellmath__48_I194 (.Y(N264), .A(N196), .B(N212), .S0(N540));
MXI2XL inst_cellmath__48_I195 (.Y(N265), .A(N197), .B(N213), .S0(N540));
MXI2XL inst_cellmath__48_I196 (.Y(N266), .A(N198), .B(N214), .S0(N540));
MXI2XL inst_cellmath__48_I197 (.Y(N267), .A(N199), .B(N215), .S0(N540));
MXI2XL inst_cellmath__48_I198 (.Y(N268), .A(N200), .B(N216), .S0(N540));
MXI2XL inst_cellmath__48_I199 (.Y(N269), .A(N201), .B(N217), .S0(N538));
MXI2XL inst_cellmath__48_I200 (.Y(N270), .A(N202), .B(N218), .S0(N538));
MXI2XL inst_cellmath__48_I201 (.Y(N271), .A(N203), .B(N219), .S0(N538));
MXI2X1 inst_cellmath__48_I202 (.Y(N272), .A(N204), .B(N220), .S0(N538));
MXI2X1 inst_cellmath__48_I203 (.Y(N273), .A(N205), .B(N221), .S0(N538));
MXI2X1 inst_cellmath__48_I204 (.Y(N274), .A(N206), .B(N222), .S0(N537));
MXI2XL inst_cellmath__48_I205 (.Y(N275), .A(N207), .B(N224), .S0(N537));
MXI2XL inst_cellmath__48_I206 (.Y(N276), .A(N208), .B(N226), .S0(N537));
MXI2XL inst_cellmath__48_I207 (.Y(N277), .A(N209), .B(N228), .S0(N537));
NOR2XL inst_cellmath__48_I208 (.Y(N278), .A(N210), .B(N537));
NOR2XL inst_cellmath__48_I209 (.Y(N280), .A(N211), .B(N536));
NOR2XL inst_cellmath__48_I210 (.Y(N282), .A(N212), .B(N536));
NOR2XL inst_cellmath__48_I211 (.Y(N284), .A(N213), .B(N536));
NOR2XL inst_cellmath__48_I212 (.Y(N286), .A(N214), .B(N536));
NOR2XL inst_cellmath__48_I213 (.Y(N288), .A(N215), .B(N536));
NOR2XL inst_cellmath__48_I214 (.Y(N290), .A(N216), .B(N535));
NOR2XL inst_cellmath__48_I215 (.Y(N292), .A(N217), .B(N535));
NOR2XL inst_cellmath__48_I216 (.Y(N294), .A(N218), .B(N535));
NOR2X1 inst_cellmath__48_I217 (.Y(N296), .A(N219), .B(N535));
NOR2XL inst_cellmath__48_I218 (.Y(N298), .A(N220), .B(N535));
NOR2XL inst_cellmath__48_I219 (.Y(N300), .A(N221), .B(N534));
NOR2XL inst_cellmath__48_I220 (.Y(N302), .A(N222), .B(N534));
NOR2XL inst_cellmath__48_I221 (.Y(N304), .A(N224), .B(N534));
NOR2XL inst_cellmath__48_I222 (.Y(N306), .A(N226), .B(N534));
NOR2XL inst_cellmath__48_I223 (.Y(N308), .A(N228), .B(N534));
INVXL inst_cellmath__48_I417 (.Y(N541), .A(inst_cellmath__48_in0[3]));
INVXL inst_cellmath__48_I418 (.Y(N542), .A(N541));
INVXL inst_cellmath__48_I423 (.Y(N547), .A(N542));
INVXL inst_cellmath__48_I422 (.Y(N546), .A(N542));
INVXL inst_cellmath__48_I421 (.Y(N545), .A(N542));
INVXL inst_cellmath__48_I420 (.Y(N544), .A(N542));
INVXL inst_cellmath__48_I419 (.Y(N543), .A(N542));
MXI2XL inst_cellmath__48_I258 (.Y(N344), .A(N272), .B(N264), .S0(N547));
MXI2XL inst_cellmath__48_I259 (.Y(N345), .A(N273), .B(N265), .S0(N547));
MXI2XL inst_cellmath__48_I260 (.Y(N346), .A(N274), .B(N266), .S0(N547));
MXI2XL inst_cellmath__48_I261 (.Y(N347), .A(N275), .B(N267), .S0(N547));
MXI2XL inst_cellmath__48_I262 (.Y(N348), .A(N276), .B(N268), .S0(N547));
MXI2X1 inst_cellmath__48_I263 (.Y(N349), .A(N277), .B(N269), .S0(N546));
MXI2X1 inst_cellmath__48_I264 (.Y(N350), .A(N278), .B(N270), .S0(N546));
MXI2XL inst_cellmath__48_I265 (.Y(N351), .A(N280), .B(N271), .S0(N546));
MXI2X1 inst_cellmath__48_I266 (.Y(N352), .A(N282), .B(N272), .S0(N546));
MXI2X1 inst_cellmath__48_I267 (.Y(N353), .A(N284), .B(N273), .S0(N546));
MXI2X1 inst_cellmath__48_I268 (.Y(N354), .A(N286), .B(N274), .S0(N545));
MXI2X1 inst_cellmath__48_I269 (.Y(N355), .A(N288), .B(N275), .S0(N545));
MXI2XL inst_cellmath__48_I270 (.Y(N356), .A(N290), .B(N276), .S0(N545));
MXI2XL inst_cellmath__48_I271 (.Y(N357), .A(N292), .B(N277), .S0(N545));
MXI2XL inst_cellmath__48_I272 (.Y(N358), .A(N294), .B(N278), .S0(N545));
MXI2XL inst_cellmath__48_I273 (.Y(N359), .A(N296), .B(N280), .S0(N544));
MXI2XL inst_cellmath__48_I274 (.Y(N360), .A(N298), .B(N282), .S0(N544));
MXI2XL inst_cellmath__48_I275 (.Y(N361), .A(N300), .B(N284), .S0(N544));
MXI2XL inst_cellmath__48_I276 (.Y(N362), .A(N302), .B(N286), .S0(N544));
MXI2XL inst_cellmath__48_I277 (.Y(N363), .A(N304), .B(N288), .S0(N544));
MXI2XL inst_cellmath__48_I278 (.Y(N364), .A(N306), .B(N290), .S0(N543));
MXI2XL inst_cellmath__48_I279 (.Y(N365), .A(N308), .B(N292), .S0(N543));
NAND2XL inst_cellmath__48_I280 (.Y(N366), .A(N294), .B(N543));
NAND2X2 inst_cellmath__48_I281 (.Y(N368), .A(N296), .B(N543));
NAND2XL inst_cellmath__48_I282 (.Y(N370), .A(N298), .B(N543));
INVXL inst_cellmath__48_I424 (.Y(N548), .A(inst_cellmath__48_in0[5]));
INVXL inst_cellmath__48_I425 (.Y(N549), .A(N548));
INVXL inst_cellmath__48_I426 (.Y(N550), .A(N549));
INVXL inst_cellmath__48_I431 (.Y(N555), .A(N550));
INVXL inst_cellmath__48_I430 (.Y(N554), .A(N550));
INVXL inst_cellmath__48_I429 (.Y(N553), .A(N550));
INVXL inst_cellmath__48_I428 (.Y(N552), .A(N550));
INVXL inst_cellmath__48_I427 (.Y(N551), .A(N550));
NOR2XL inst_cellmath__48_I322 (.Y(inst_cellmath__48_out0[0]), .A(N344), .B(N555));
NOR2XL inst_cellmath__48_I323 (.Y(inst_cellmath__48_out0[1]), .A(N345), .B(N555));
NOR2X1 inst_cellmath__48_I324 (.Y(inst_cellmath__48_out0[2]), .A(N346), .B(N555));
NOR2XL inst_cellmath__48_I325 (.Y(inst_cellmath__48_out0[3]), .A(N347), .B(N555));
NOR2XL inst_cellmath__48_I326 (.Y(inst_cellmath__48_out0[4]), .A(N348), .B(N555));
NOR2X1 inst_cellmath__48_I327 (.Y(inst_cellmath__48_out0[5]), .A(N349), .B(N554));
NOR2X1 inst_cellmath__48_I328 (.Y(inst_cellmath__48_out0[6]), .A(N350), .B(N554));
NOR2XL inst_cellmath__48_I329 (.Y(inst_cellmath__48_out0[7]), .A(N351), .B(N554));
NOR2X2 inst_cellmath__48_I330 (.Y(inst_cellmath__48_out0[8]), .A(N352), .B(N554));
NOR2X1 inst_cellmath__48_I331 (.Y(inst_cellmath__48_out0[9]), .A(N353), .B(N554));
NOR2X1 inst_cellmath__48_I332 (.Y(inst_cellmath__48_out0[10]), .A(N354), .B(N553));
NOR2X1 inst_cellmath__48_I333 (.Y(inst_cellmath__48_out0[11]), .A(N355), .B(N553));
NOR2XL inst_cellmath__48_I334 (.Y(inst_cellmath__48_out0[12]), .A(N356), .B(N553));
NOR2XL inst_cellmath__48_I335 (.Y(inst_cellmath__48_out0[13]), .A(N357), .B(N553));
NOR2XL inst_cellmath__48_I336 (.Y(inst_cellmath__48_out0[14]), .A(N358), .B(N553));
NOR2XL inst_cellmath__48_I337 (.Y(inst_cellmath__48_out0[15]), .A(N359), .B(N552));
NOR2XL inst_cellmath__48_I338 (.Y(inst_cellmath__48_out0[16]), .A(N360), .B(N552));
NOR2XL inst_cellmath__48_I339 (.Y(inst_cellmath__48_out0[17]), .A(N361), .B(N552));
NOR2XL inst_cellmath__48_I340 (.Y(inst_cellmath__48_out0[18]), .A(N362), .B(N552));
NOR2XL inst_cellmath__48_I341 (.Y(inst_cellmath__48_out0[19]), .A(N363), .B(N552));
NOR2XL inst_cellmath__48_I342 (.Y(inst_cellmath__48_out0[20]), .A(N364), .B(N551));
NOR2XL inst_cellmath__48_I343 (.Y(inst_cellmath__48_out0[21]), .A(N365), .B(N551));
NOR2XL inst_cellmath__48_I344 (.Y(inst_cellmath__48_out0[22]), .A(N366), .B(N551));
NOR2X4 inst_cellmath__48_I345 (.Y(inst_cellmath__48_out0[23]), .A(N368), .B(N551));
NOR2XL inst_cellmath__48_I346 (.Y(inst_cellmath__48_out0[24]), .A(N370), .B(N551));
endmodule

module cynw_cm_float_sin_inst_cellmath__61_0_bdw1946085813_bdw (
	inst_cellmath__61_0_out0,
	inst_cellmath__61_0_in0
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__61_0_out0;
input [23:0] inst_cellmath__61_0_in0;
wire N100,N163,N164;
INVXL inst_cellmath__61_0_I51 (.Y(N100), .A(inst_cellmath__61_0_in0[5]));
CLKINVX6 inst_cellmath__61_0_I109 (.Y(N163), .A(inst_cellmath__61_0_in0[23]));
CLKINVX8 inst_cellmath__61_0_I110 (.Y(N164), .A(N163));
XOR2XL inst_cellmath__61_0_I320 (.Y(inst_cellmath__61_0_out0[0]), .A(inst_cellmath__61_0_in0[0]), .B(N164));
XOR2XL inst_cellmath__61_0_I321 (.Y(inst_cellmath__61_0_out0[1]), .A(inst_cellmath__61_0_in0[1]), .B(N164));
XOR2XL inst_cellmath__61_0_I322 (.Y(inst_cellmath__61_0_out0[2]), .A(inst_cellmath__61_0_in0[2]), .B(N164));
XOR2XL inst_cellmath__61_0_I323 (.Y(inst_cellmath__61_0_out0[3]), .A(inst_cellmath__61_0_in0[3]), .B(N164));
XOR2XL inst_cellmath__61_0_I324 (.Y(inst_cellmath__61_0_out0[4]), .A(inst_cellmath__61_0_in0[4]), .B(N164));
MXI2X1 inst_cellmath__61_0_I74 (.Y(inst_cellmath__61_0_out0[5]), .A(N100), .B(inst_cellmath__61_0_in0[5]), .S0(N164));
XOR2XL inst_cellmath__61_0_I326 (.Y(inst_cellmath__61_0_out0[6]), .A(inst_cellmath__61_0_in0[6]), .B(N164));
XOR2XL inst_cellmath__61_0_I327 (.Y(inst_cellmath__61_0_out0[7]), .A(inst_cellmath__61_0_in0[7]), .B(N164));
XOR2XL inst_cellmath__61_0_I328 (.Y(inst_cellmath__61_0_out0[8]), .A(inst_cellmath__61_0_in0[8]), .B(N164));
XOR2XL inst_cellmath__61_0_I201 (.Y(inst_cellmath__61_0_out0[9]), .A(inst_cellmath__61_0_in0[9]), .B(N164));
XOR2XL inst_cellmath__61_0_I329 (.Y(inst_cellmath__61_0_out0[10]), .A(inst_cellmath__61_0_in0[10]), .B(N164));
XOR2XL inst_cellmath__61_0_I330 (.Y(inst_cellmath__61_0_out0[11]), .A(inst_cellmath__61_0_in0[11]), .B(N164));
XOR2XL inst_cellmath__61_0_I331 (.Y(inst_cellmath__61_0_out0[12]), .A(inst_cellmath__61_0_in0[12]), .B(N164));
XOR2XL inst_cellmath__61_0_I332 (.Y(inst_cellmath__61_0_out0[13]), .A(inst_cellmath__61_0_in0[13]), .B(N164));
XOR2XL inst_cellmath__61_0_I333 (.Y(inst_cellmath__61_0_out0[14]), .A(inst_cellmath__61_0_in0[14]), .B(N164));
XOR2XL inst_cellmath__61_0_I138 (.Y(inst_cellmath__61_0_out0[15]), .A(inst_cellmath__61_0_in0[15]), .B(N164));
XOR2XL inst_cellmath__61_0_I334 (.Y(inst_cellmath__61_0_out0[16]), .A(inst_cellmath__61_0_in0[16]), .B(N164));
XOR2XL inst_cellmath__61_0_I140 (.Y(inst_cellmath__61_0_out0[17]), .A(inst_cellmath__61_0_in0[17]), .B(N164));
XOR2XL inst_cellmath__61_0_I141 (.Y(inst_cellmath__61_0_out0[18]), .A(inst_cellmath__61_0_in0[18]), .B(N164));
XOR2XL inst_cellmath__61_0_I142 (.Y(inst_cellmath__61_0_out0[19]), .A(inst_cellmath__61_0_in0[19]), .B(N164));
XOR2XL inst_cellmath__61_0_I143 (.Y(inst_cellmath__61_0_out0[20]), .A(inst_cellmath__61_0_in0[20]), .B(N164));
XOR2XL inst_cellmath__61_0_I144 (.Y(inst_cellmath__61_0_out0[21]), .A(inst_cellmath__61_0_in0[21]), .B(N164));
XOR2XL inst_cellmath__61_0_I145 (.Y(inst_cellmath__61_0_out0[22]), .A(inst_cellmath__61_0_in0[22]), .B(N164));
endmodule

module cynw_cm_float_sin_inst_cellmath__195__80__2WWMM_2WWMM_bdw1946085813_bdw (
	inst_cellmath__195__80__2WWMM_2WWMM_out0,
	inst_cellmath__195__80__2WWMM_2WWMM_in0
	); /* architecture "gate_level" */ 
output [72:0] inst_cellmath__195__80__2WWMM_2WWMM_out0;
input [22:17] inst_cellmath__195__80__2WWMM_2WWMM_in0;
wire N82,N85,N88,N89,N91,N92,N93 
	,N95,N96,N98,N102,N104,N106,N107,N108 
	,N110,N111,N112,N113,N114,N116,N117,N118 
	,N119,N122,N123,N124,N126,N128,N129,N131 
	,N133,N134,N135,N136,N137,N138,N141,N142 
	,N143,N144,N145,N146,N147,N149,N150,N151 
	,N152,N153,N154,N155,N156,N159,N160,N161 
	,N163,N164,N167,N168,N169,N170,N173,N174 
	,N4258,N4260,N4261,N4262,N4263,N4267,N4268,N4272 
	,N4273,N4274,N4276,N4277,N4278,N4280,N4281,N4288 
	,N4289,N4290,N4291,N4292,N4293,N4294,N4296,N4297 
	,N4298,N4302,N4303,N4304,N4305,N4307,N4309,N4310 
	,N4319,N4321,N4322,N4323,N4324,N4325,N4326,N4327 
	,N4329,N4330,N4331,N4332,N4333,N4336,N4337,N4338 
	,N4339,N4347,N4348,N4350,N4351,N4358,N4361,N4362 
	,N4363,N4364,N4365,N4366,N4367,N4368,N4370,N4371 
	,N4384,N4389,N4393,N4396,N4400,N4401,N4410,N4413 
	,N4415,N4416,N4419,N4421,N4422,N4425,N4428,N4429 
	,N4436,N4438,N4442,N4443,N4444,N4446,N4448,N4449 
	,N4451,N4452,N4454,N4455,N4456,N4459,N4460,N4462 
	,N4471,N4475,N4477,N4480,N4481,N4484,N4485,N4486 
	,N4488,N4490,N4491,N4493,N4494,N4500,N4503,N4507 
	,N4511,N4514,N4515,N4516,N4517,N4521,N4522,N4527 
	,N4528,N4534,N4535,N4537,N4538,N4539,N4541,N4542 
	,N4548,N4549,N4550,N4552,N4553,N4554,N4555,N4556 
	,N4560,N4561,N4562,N4574,N4575,N4576,N4585,N4586 
	,N4587,N4588,N4589,N4590,N4591,N4594,N4597,N4603 
	,N4607,N4608,N4609,N4610,N4614,N4618,N4621,N4625 
	,N4627,N4628,N4631,N4634,N4635,N4643,N4645,N4647 
	,N4652,N4654,N4656,N4659,N4661,N4667,N4668,N4669 
	,N4677,N4678,N4682,N4684,N4685,N4686,N4688,N4689 
	,N4692,N4696,N4697,N4699,N4702,N4704,N4706,N4707 
	,N4708,N4710,N4718,N4719,N4723,N4724,N4731,N4732 
	,N4733,N4735,N4736,N4737,N4740,N4741,N4743,N4744 
	,N4755,N4762,N4765,N4767,N4769,N4771,N4772,N4773 
	,N4774,N4778,N4784,N4789,N4790,N4794,N4795,N4799 
	,N4801,N4802,N4804,N4805,N4807,N4809,N4810,N4821 
	,N4822,N4824,N4825,N4826,N4827,N4829,N4831,N4832 
	,N4835,N4839,N4842,N4846,N4847,N4860,N4865,N4866 
	,N4875,N4876,N4886,N4887,N4893,N4897,N4900,N4901 
	,N4902,N4915,N4917,N4919,N4922,N4924,N4937,N4940 
	,N4943,N4945,N4946,N4948,N4950,N4952,N4953,N4979 
	,N4980,N4984,N4991,N4992,N4993,N4995,N4998,N5002 
	,N5005,N5014,N5017,N5019,N5020,N5025,N5031,N5035 
	,N5036,N5038,N5055,N5056,N5061,N5063,N5065,N5067 
	,N5069,N5078,N5081,N5090,N5096,N5098,N5099,N5102 
	,N5110,N5116,N5126,N5127,N5128,N5129,N5131,N5134 
	,N5135,N5136,N5139,N5140,N5148,N5155,N5156,N5161 
	,N5163,N5164,N5167,N5168,N5170,N5172,N5184,N5185 
	,N5190,N5198,N5201,N5203,N5204,N5205,N5218,N5223 
	,N5224,N5225,N5226,N5229,N5230,N5236,N5238,N5240 
	,N5243,N5260,N5261,N5263,N5264,N5265,N5267,N5270 
	,N5272,N5273,N5285,N5287,N5294,N5298,N5300,N5302 
	,N5304,N5306,N5308,N5311,N5321,N5324,N5330,N5331 
	,N5335,N5339,N5340,N5342,N5350,N5353,N5355,N5358 
	,N5363,N5366,N5368,N5369,N5370,N5371,N5374,N5375 
	,N5376,N5385,N5394,N5396,N5399,N5402,N5406,N5410 
	,N5420,N5423,N5427,N5429,N5435,N5438,N5439,N5442 
	,N5447,N5454,N5461,N5465,N5466,N5467,N5474,N5481 
	,N5482,N5485,N5486,N5497,N5498,N5505,N5507,N5508 
	,N5512,N5517,N5518,N5539,N5544,N5545,N5547,N5560 
	,N5562,N5566,N5570,N5572,N5574,N5575,N5576,N5579 
	,N5582,N5583,N5593,N5594,N5595,N5596,N5604,N5608 
	,N5609,N5610,N5613,N5614,N5635,N5639,N5641,N5642 
	,N5643,N5654,N5657,N5662,N5664,N5669,N5671,N5675 
	,N5680,N5682,N5689,N5694,N5702,N5707,N5708,N5713 
	,N5714,N5731,N5738,N5741,N5742,N5744,N5746,N5748 
	,N5751,N5768,N5771,N5772,N5773,N5774,N5777,N5779 
	,N5781,N5791,N5801,N5803,N5804,N5805,N5806,N5808 
	,N5809,N5812,N5821,N5823,N5835,N5838,N5839,N5842 
	,N5853,N5861,N5864,N5865,N5866,N5869,N5872,N5874 
	,N5875,N5884,N5885,N5886,N5892,N5900,N5903,N5906 
	,N5908,N5910,N5919,N5927,N5928,N5930,N5935,N5936 
	,N5938,N5939,N5942,N5943,N5963,N5967,N5970,N5971 
	,N5974,N5975,N5977,N5996,N5998,N6004,N6006,N6010 
	,N6011,N6023,N6025,N6032,N6034,N6036,N6038,N6049 
	,N6055,N6062,N6065,N6067,N6068,N6070,N6072,N6073 
	,N6074,N6086,N6096,N6101,N6102,N6104,N6109,N6110 
	,N6113,N6114,N6121,N6129,N6135,N6138,N6139,N6142 
	,N6144,N6145,N6147,N6149,N6160,N6172,N6174,N6175 
	,N6178,N6181,N6183,N6187,N6189,N6195,N6207,N6212 
	,N6213,N6214,N6216,N6218,N6220,N6230,N6231,N6245 
	,N6247,N6251,N6263,N6264,N6267,N6272,N6277,N6278 
	,N6279,N6280,N6287,N6298,N6301,N6303,N6312,N6313 
	,N6314,N6315,N6316,N6317,N6320,N6323,N6344,N6345 
	,N6346,N6350,N6354,N6356,N6358,N6361,N6362,N6364 
	,N6383,N6389,N6391,N6395,N6396,N6397,N6418,N6420 
	,N6422,N6426,N6429,N6432,N6435,N6447,N6453,N6457 
	,N6459,N6461,N6463,N6465,N6466,N6467,N6485,N6495 
	,N6497,N6500,N6501,N6502,N6503,N6508,N6509,N6511 
	,N6517,N6523,N6525,N6531,N6536,N6539,N6549,N6558 
	,N6563,N6564,N6568,N6569,N6570,N6591,N6592,N6593 
	,N6594,N6595,N6601,N6624,N6625,N6626,N6631,N6632 
	,N6633,N6640,N6654,N6656,N6658,N6660,N6669,N6675 
	,N6679,N6685,N6689,N6695,N6697,N6701,N6705,N6707 
	,N6711,N6713,N6715,N6719,N6721,N6727,N6733,N6739 
	,N6743,N6753,N6755,N6769,N6777,N6787,N6789,N6791 
	,N6793,N6795,N6797,N6799,N6801,N6805,N6807,N6809 
	,N6811,N6813,N6815,N6817,N6823,N6833,N6835,N6837 
	,N8068,N8071,N8072,N8073,N8076,N8079,N8080,N8081 
	,N8090,N8091,N8092,N8095,N8096,N8097,N8098,N8099 
	,N8100,N8103,N8106,N8107,N8108,N8109,N8110,N8111 
	,N8112,N8113,N8114,N8117,N8118,N8119,N8126,N8127 
	,N8128,N8129,N8130,N8137,N8138,N8139,N8142,N8143 
	,N8144,N8150,N8151,N8152,N8161,N8162,N8163,N8168 
	,N8174,N8175,N8176,N8178,N8182,N8185,N8186,N8187 
	,N8188,N8189,N8198,N8202,N8206,N8210,N8211,N8212 
	,N8213,N8216,N8218,N8219,N8223,N8227,N8233,N8234 
	,N8238,N8242,N8247,N8248,N8249,N8250,N8255,N8256 
	,N8257,N8259,N8260,N8264,N8277,N8281,N8284,N8288 
	,N8294,N8299,N8304,N8308,N8309,N8310,N8311,N8315 
	,N8319,N8322,N8324,N8325,N8332,N8336,N8339,N8346 
	,N8350,N8354,N8362,N8366,N8371,N8372,N8375,N8379 
	,N8383,N8386,N8388,N8390,N8394,N8397,N8401,N8402 
	,N8407,N8411,N8413,N8417,N8421,N8426,N8427,N8428 
	,N8429,N8430,N8435,N8439,N8442,N8444,N8445,N8449 
	,N8455,N8459,N8460,N8461,N8462,N8464,N8467,N8470 
	,N8474,N8478,N8479,N8481,N8482,N8486,N8487,N8496 
	,N8500,N8505,N8506,N8508,N8509,N8512,N8513,N8514 
	,N8515,N8521,N8525,N8528,N8529,N8535,N8539,N8543 
	,N8544,N8546,N8547,N8551,N8562,N8567,N8575,N8579 
	,N8594,N8595,N8598,N8601,N8602,N8603,N8605,N8607 
	,N8609,N8621,N8628,N8635,N8644,N8650,N8657,N8664 
	,N8671,N8678,N8685,N8692,N8699,N8706,N8713,N8722 
	,N8728,N8735,N8742,N8749,N8756,N8763,N8770,N8779 
	,N8787,N8793,N8800,N8807,N8816,N8824,N8832,N8838 
	,N8847,N8855,N8863,N8869,N8876,N8885,N8893,N8901 
	,N8907,N8914,N8921,N8928,N8937,N8943,N8952,N8960 
	,N8966,N8973,N8982,N8988,N8997,N9003,N9010,N9017 
	,N9026,N9032,N9039,N9048,N9056,N9064,N9070,N9077 
	,N11605,N11613,N11621;
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5007 (.Y(N8068), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1 (.Y(N82), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I7095 (.Y(N8071), .A(N82), .B(N8068));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5012 (.Y(N8073), .A(N8071));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5011 (.Y(N8072), .A(N8071));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5015 (.Y(N8076), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4 (.Y(N85), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I7227 (.Y(N8079), .A(N85), .B(N8076));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5020 (.Y(N8081), .A(N8079));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5019 (.Y(N8080), .A(N8079));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I6 (.Y(N6669), .A(N8081), .B(N8073));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I7 (.Y(N88), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I8 (.Y(N89), .A(N88), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10033 (.Y(N8090), .A(N8076), .B(N89));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5031 (.Y(N8092), .A(N8090));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5030 (.Y(N8091), .A(N8090));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10 (.Y(N91), .A(N8092), .B(N8073));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I11 (.Y(N92), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[18]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I12 (.Y(N93), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[17]), .B(N92));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I7099 (.Y(N8095), .A(N8076), .B(N93));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5036 (.Y(N8097), .A(N8095));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5035 (.Y(N8096), .A(N8095));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I14 (.Y(N95), .A(N8097), .B(N8073));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I15 (.Y(N96), .A(N88), .B(N92));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I16 (.Y(N6675), .A(N96), .B(N8076));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5037 (.Y(N8098), .A(N6675));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5039 (.Y(N8100), .A(N8098));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5038 (.Y(N8099), .A(N8098));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I17 (.Y(N98), .A(N8100), .B(N8072));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10035 (.Y(N8103), .A(N85), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I19 (.Y(N6679), .A(N8103), .B(N8072));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I5650 (.Y(N8106), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]), .B(N89));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5047 (.Y(N8108), .A(N8106));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5046 (.Y(N8107), .A(N8106));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I21 (.Y(N102), .A(N8108), .B(N8072));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10036 (.Y(N8109), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]), .B(N93));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5050 (.Y(N8111), .A(N8109));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5049 (.Y(N8110), .A(N8109));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I23 (.Y(N104), .A(N8111), .B(N8072));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I24 (.Y(N6685), .A(N96), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[19]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I5051 (.Y(N8112), .A(N6685));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5053 (.Y(N8114), .A(N8112));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5052 (.Y(N8113), .A(N8112));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I25 (.Y(N106), .A(N8114), .B(N8072));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I26 (.Y(N107), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I27 (.Y(N108), .A(N107), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10038 (.Y(N8117), .A(N8068), .B(N108));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5058 (.Y(N8119), .A(N8117));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5057 (.Y(N8118), .A(N8117));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I29 (.Y(N110), .A(N8081), .B(N8119));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I30 (.Y(N111), .A(N8092), .B(N8119));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I31 (.Y(N112), .A(N8097), .B(N8119));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I32 (.Y(N113), .A(N8100), .B(N8118));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I33 (.Y(N114), .A(N8103), .B(N8118));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I34 (.Y(N6689), .A(N8108), .B(N8118));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I35 (.Y(N116), .A(N8111), .B(N8118));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I36 (.Y(N117), .A(N8114), .B(N8118));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I37 (.Y(N118), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[21]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I38 (.Y(N119), .A(inst_cellmath__195__80__2WWMM_2WWMM_in0[20]), .B(N118));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10039 (.Y(N8126), .A(N119), .B(N8068));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5067 (.Y(N8128), .A(N8126));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5066 (.Y(N8127), .A(N8126));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10040 (.Y(N8129), .A(N8081), .B(N8128));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5069 (.Y(N8130), .A(N8129));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I41 (.Y(N122), .A(N8092), .B(N8128));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I42 (.Y(N123), .A(N8097), .B(N8128));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I43 (.Y(N124), .A(N8100), .B(N8127));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I44 (.Y(N6695), .A(N8103), .B(N8127));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I45 (.Y(N126), .A(N8108), .B(N8127));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I46 (.Y(N6697), .A(N8111), .B(N8127));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I47 (.Y(N128), .A(N8114), .B(N8127));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I48 (.Y(N129), .A(N107), .B(N118));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I7107 (.Y(N8137), .A(N129), .B(N8068));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5078 (.Y(N8139), .A(N8137));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5077 (.Y(N8138), .A(N8137));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I50 (.Y(N131), .A(N8080), .B(N8139));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I51 (.Y(N6701), .A(N8091), .B(N8139));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I52 (.Y(N133), .A(N8096), .B(N8139));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I53 (.Y(N134), .A(N8099), .B(N8138));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I54 (.Y(N135), .A(N8103), .B(N8138));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I55 (.Y(N136), .A(N8107), .B(N8138));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I56 (.Y(N137), .A(N8110), .B(N8138));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I57 (.Y(N138), .A(N8113), .B(N8138));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10041 (.Y(N8142), .A(N82), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5083 (.Y(N8144), .A(N8142));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5082 (.Y(N8143), .A(N8142));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I59 (.Y(N6705), .A(N8080), .B(N8144));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I60 (.Y(N141), .A(N8091), .B(N8144));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I61 (.Y(N142), .A(N8096), .B(N8144));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I62 (.Y(N143), .A(N8099), .B(N8143));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I63 (.Y(N144), .A(N8103), .B(N8143));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I64 (.Y(N145), .A(N8107), .B(N8143));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I65 (.Y(N146), .A(N8110), .B(N8143));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I66 (.Y(N147), .A(N8113), .B(N8143));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I67 (.Y(N6707), .A(N108), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I68 (.Y(N149), .A(N8080), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I69 (.Y(N150), .A(N8091), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I70 (.Y(N151), .A(N8096), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I71 (.Y(N152), .A(N8099), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I72 (.Y(N153), .A(N8103), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I73 (.Y(N154), .A(N8107), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I74 (.Y(N155), .A(N8110), .B(N6707));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I75 (.Y(N156), .A(N8113), .B(N6707));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10042 (.Y(N8150), .A(N119), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5091 (.Y(N8152), .A(N8150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5090 (.Y(N8151), .A(N8150));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I77 (.Y(N6711), .A(N8080), .B(N8152));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I78 (.Y(N159), .A(N8091), .B(N8152));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I79 (.Y(N160), .A(N8096), .B(N8152));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I80 (.Y(N161), .A(N8099), .B(N8151));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I81 (.Y(N6713), .A(N8103), .B(N8151));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I82 (.Y(N163), .A(N8107), .B(N8151));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I83 (.Y(N164), .A(N8110), .B(N8151));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I84 (.Y(N6715), .A(N8113), .B(N8151));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10043 (.Y(N8161), .A(N129), .B(inst_cellmath__195__80__2WWMM_2WWMM_in0[22]));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5102 (.Y(N8163), .A(N8161));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5101 (.Y(N8162), .A(N8161));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I86 (.Y(N167), .A(N8080), .B(N8163));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I87 (.Y(N168), .A(N8091), .B(N8163));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I88 (.Y(N169), .A(N8096), .B(N8163));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I89 (.Y(N170), .A(N8099), .B(N8162));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I90 (.Y(N6719), .A(N8103), .B(N8162));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I91 (.Y(N6721), .A(N8107), .B(N8162));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I92 (.Y(N173), .A(N8110), .B(N8162));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I93 (.Y(N174), .A(N8113), .B(N8162));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5107 (.Y(N8168), .A(N6669));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5113 (.Y(N8174), .A(N91));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5662 (.Y(N8175), .A(N91), .B(N6669));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5117 (.Y(N8178), .A(N8175));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5115 (.Y(N8176), .A(N8175));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5121 (.Y(N8182), .A(N95));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5125 (.Y(N8186), .A(N98));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5124 (.Y(N8185), .A(N98));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7112 (.Y(N8187), .A(N98), .B(N95));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5128 (.Y(N8189), .A(N8187));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5127 (.Y(N8188), .A(N8187));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I249 (.Y(N6727), .A(N102), .B(N6679));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5137 (.Y(N8198), .A(N102));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5141 (.Y(N8202), .A(N6679));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5145 (.Y(N8206), .A(N104));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5149 (.Y(N8210), .A(N106));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7114 (.Y(N8211), .A(N106), .B(N104));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5152 (.Y(N8213), .A(N8211));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5151 (.Y(N8212), .A(N8211));
OR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10044 (.Y(N8216), .A(N111), .B(N110));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5158 (.Y(N8219), .A(N8216));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5157 (.Y(N8218), .A(N8216));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5162 (.Y(N8223), .A(N110));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5166 (.Y(N8227), .A(N111));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I477 (.Y(N6733), .A(N113), .B(N112));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5173 (.Y(N8234), .A(N113));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5172 (.Y(N8233), .A(N113));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5177 (.Y(N8238), .A(N112));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5181 (.Y(N8242), .A(N6689));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5186 (.Y(N8247), .A(N114));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5678 (.Y(N8248), .A(N6689), .B(N114));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5189 (.Y(N8250), .A(N8248));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5188 (.Y(N8249), .A(N8248));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5195 (.Y(N8256), .A(N116));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5194 (.Y(N8255), .A(N116));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10045 (.Y(N8257), .A(N117), .B(N116));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5199 (.Y(N8260), .A(N8257));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5198 (.Y(N8259), .A(N8257));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5203 (.Y(N8264), .A(N117));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I707 (.Y(N6739), .A(N122), .B(N8130));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5216 (.Y(N8277), .A(N122));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5220 (.Y(N8281), .A(N124));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10046 (.Y(N8284), .A(N124), .B(N123));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5227 (.Y(N8288), .A(N123));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I857 (.Y(N6743), .A(N126), .B(N6695));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5233 (.Y(N8294), .A(N6695));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5238 (.Y(N8299), .A(N126));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5243 (.Y(N8304), .A(N128));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5247 (.Y(N8308), .A(N6697));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7123 (.Y(N8309), .A(N128), .B(N6697));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5250 (.Y(N8311), .A(N8309));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5249 (.Y(N8310), .A(N8309));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5254 (.Y(N8315), .A(N6701));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5258 (.Y(N8319), .A(N131));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10047 (.Y(N8322), .A(N6701), .B(N131));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5264 (.Y(N8325), .A(N8322));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5263 (.Y(N8324), .A(N8322));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5271 (.Y(N8332), .A(N134));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10048 (.Y(N8336), .A(N134), .B(N133));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5278 (.Y(N8339), .A(N133));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10049 (.Y(N8346), .A(N136), .B(N135));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5289 (.Y(N8350), .A(N136));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5293 (.Y(N8354), .A(N135));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1237 (.Y(N6753), .A(N138), .B(N137));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5301 (.Y(N8362), .A(N137));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5305 (.Y(N8366), .A(N138));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1313 (.Y(N6755), .A(N141), .B(N6705));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5310 (.Y(N8371), .A(N6705));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5311 (.Y(N8372), .A(N141));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5314 (.Y(N8375), .A(N143));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5318 (.Y(N8379), .A(N142));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10050 (.Y(N8383), .A(N143), .B(N142));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5325 (.Y(N8386), .A(N144));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7129 (.Y(N8388), .A(N145), .B(N144));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5329 (.Y(N8390), .A(N8388));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5333 (.Y(N8394), .A(N145));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10052 (.Y(N8397), .A(N147), .B(N146));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5341 (.Y(N8402), .A(N147));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5340 (.Y(N8401), .A(N147));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5346 (.Y(N8407), .A(N146));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5350 (.Y(N8411), .A(N149));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I7250 (.Y(N8413), .A(N150), .B(N149));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5356 (.Y(N8417), .A(N150));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5360 (.Y(N8421), .A(N152));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5366 (.Y(N8427), .A(N151));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5365 (.Y(N8426), .A(N151));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7132 (.Y(N8428), .A(N152), .B(N151));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5369 (.Y(N8430), .A(N8428));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5368 (.Y(N8429), .A(N8428));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5374 (.Y(N8435), .A(N153));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5378 (.Y(N8439), .A(N154));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10053 (.Y(N8442), .A(N154), .B(N153));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5384 (.Y(N8445), .A(N8442));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5383 (.Y(N8444), .A(N8442));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5388 (.Y(N8449), .A(N156));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1852 (.Y(N6769), .A(N156), .B(N155));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5394 (.Y(N8455), .A(N155));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5399 (.Y(N8460), .A(N159));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5398 (.Y(N8459), .A(N159));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I7252 (.Y(N8461), .A(N159), .B(N6711));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5403 (.Y(N8464), .A(N8461));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5401 (.Y(N8462), .A(N8461));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5406 (.Y(N8467), .A(N6711));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10054 (.Y(N8470), .A(N161), .B(N160));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5413 (.Y(N8474), .A(N161));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5417 (.Y(N8478), .A(N160));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10055 (.Y(N8479), .A(N163), .B(N6713));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I5421 (.Y(N8482), .A(N8479));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5420 (.Y(N8481), .A(N8479));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5425 (.Y(N8486), .A(N6713));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5426 (.Y(N8487), .A(N163));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2149 (.Y(N6777), .A(N6715), .B(N164));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5435 (.Y(N8496), .A(N6715));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5439 (.Y(N8500), .A(N164));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5444 (.Y(N8505), .A(N167));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I5723 (.Y(N8506), .A(N168), .B(N167));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5448 (.Y(N8509), .A(N8506));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5447 (.Y(N8508), .A(N8506));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5452 (.Y(N8513), .A(N168));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5451 (.Y(N8512), .A(N168));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10056 (.Y(N8514), .A(N170), .B(N169));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5454 (.Y(N8515), .A(N8514));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I7139 (.Y(N8521), .A(N169));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5464 (.Y(N8525), .A(N170));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5468 (.Y(N8529), .A(N6721));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5467 (.Y(N8528), .A(N6721));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10057 (.Y(N8535), .A(N6721), .B(N6719));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5478 (.Y(N8539), .A(N6719));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5482 (.Y(N8543), .A(N174));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10058 (.Y(N8544), .A(N174), .B(N173));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5486 (.Y(N8547), .A(N8544));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5485 (.Y(N8546), .A(N8544));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5490 (.Y(N8551), .A(N173));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2531 (.Y(N4258), .A(N8168), .B(N8129));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2533 (.Y(N4260), .A(N8386), .B(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2534 (.Y(N4261), .A(N8411), .B(N8529));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5731 (.Y(N4262), .AN(N152), .B(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2536 (.Y(N4263), .A(N8375), .B(N8182));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2537 (.Y(N6787), .A(N8315), .B(N8460));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2540 (.Y(N4267), .A(N134), .B(N4258));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2541 (.Y(N4268), .A(N6733), .B(N6777));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2542 (.Y(N6789), .A(N6727), .B(N6755));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5734 (.Y(N6791), .AN(N8514), .B(N8470));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2545 (.Y(N4272), .A(N4261), .B(N4262));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2546 (.Y(N4273), .A(N4263), .B(N4268));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2547 (.Y(N4274), .A(N4260), .B(N6789));
NAND2XL hyperpropagate_3_1_A_I7419 (.Y(N8621), .A(N8219), .B(N6753));
NOR2XL hyperpropagate_3_1_A_I7420 (.Y(N4276), .A(N6791), .B(N8621));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2550 (.Y(N4277), .A(N4272), .B(N4267));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2551 (.Y(N4278), .A(N4273), .B(N4274));
NAND3XL hyperpropagate_4_1_A_I10091 (.Y(N11605), .A(N8256), .B(N6743), .C(N4276));
NOR2XL hyperpropagate_4_1_A_I10092 (.Y(N4281), .A(N6787), .B(N11605));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2553 (.Y(N4280), .A(N4277), .B(N4278));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2555 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[0]), .A(N4281), .B(N4280));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2561 (.Y(N4288), .A(N8371), .B(N8129));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2562 (.Y(N4289), .A(N8294), .B(N8505));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2563 (.Y(N4290), .A(N8223), .B(N8319));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2564 (.Y(N4291), .A(N8529), .B(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2565 (.Y(N4292), .A(N8206), .B(N8439));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2566 (.Y(N4293), .A(N8421), .B(N8186));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2567 (.Y(N4294), .A(N8346), .B(N8332));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2568 (.Y(N6793), .A(N8281), .B(N8482));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2569 (.Y(N4296), .A(N8397), .B(N8413));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2570 (.Y(N4297), .A(N8260), .B(N8462));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2571 (.Y(N4298), .A(N6753));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5501 (.Y(N8562), .A(N8515));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2575 (.Y(N4302), .A(N4290), .B(N4292));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2576 (.Y(N4303), .A(N4296), .B(N4297));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2577 (.Y(N4304), .A(N6793), .B(N4291));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2578 (.Y(N4305), .A(N4294), .B(N4293));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2580 (.Y(N4307), .A(N4304), .B(N4305));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6387 (.Y(N4310), .AN(N8515), .B(N4298), .C(N4288), .D(N4289));
NAND2XL hyperpropagate_3_1_A_I7421 (.Y(N8628), .A(N4302), .B(N4303));
NOR2XL hyperpropagate_3_1_A_I7422 (.Y(N4309), .A(N4307), .B(N8628));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2584 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[1]), .A(N4310), .B(N4309));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2591 (.Y(N4319), .A(N8234), .B(N8496));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2593 (.Y(N4321), .A(N8362), .B(N8186));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2594 (.Y(N4322), .A(N8210), .B(N8535));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2595 (.Y(N4323), .A(N6743), .B(N8346));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2596 (.Y(N4324), .A(N8445), .B(N8509));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2597 (.Y(N4325), .A(N6739), .B(N8219));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2598 (.Y(N4326), .A(N8390), .B(N8413));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2599 (.Y(N4327), .A(N8325), .B(N8336));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2600 (.Y(N6795), .A(N8515), .B(N8284));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5752 (.Y(N4329), .AN(N4319), .B(N8402), .C(N8427));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2602 (.Y(N4330), .A(N4324), .B(N143));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2603 (.Y(N4331), .A(N4322), .B(N4327));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2604 (.Y(N4332), .A(N4323), .B(N4325));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2605 (.Y(N4333), .A(N4326), .B(N4321));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2607 (.Y(N4339), .A(N6795), .B(N4329));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2608 (.Y(N4336), .A(N4330), .B(N4331));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2609 (.Y(N4337), .A(N4332), .B(N4333));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2610 (.Y(N4338), .A(N4336), .B(N4337));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2612 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[2]), .A(N4339), .B(N4338));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I7164 (.Y(N4347), .AN(N126), .B(N8528));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2619 (.Y(N4348), .A(N8304), .B(N8350));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2620 (.Y(N4490), .A(N8439), .B(N8421));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2621 (.Y(N4350), .A(N8277), .B(N8496));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2622 (.Y(N4351), .A(N8198), .B(N8372));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2624 (.Y(N4993), .A(N8402), .B(N8449));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2626 (.Y(N5779), .A(N8256), .B(N8543));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5506 (.Y(N8567), .A(N8336));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2629 (.Y(N4358), .A(N8567), .B(N167));
NAND3XL hyperpropagate_4_1_A_I10093 (.Y(N11613), .A(N6733), .B(N8394), .C(N8482));
NOR2XL hyperpropagate_4_1_A_I10094 (.Y(N4361), .A(N142), .B(N11613));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2633 (.Y(N4362), .A(N4350), .B(N4993));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2634 (.Y(N4363), .A(N6787), .B(N5779));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2635 (.Y(N4364), .A(N4490), .B(N4347));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2636 (.Y(N4365), .A(N4348));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2637 (.Y(N4366), .A(N4365), .B(N4361));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2638 (.Y(N4367), .A(N4362), .B(N4358));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2639 (.Y(N4368), .A(N4363), .B(N4364));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I10061 (.Y(N4370), .A(N8562), .B(N4351), .C(N4367));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2642 (.Y(N4371), .A(N4368), .B(N4366));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2643 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[3]), .A(N4370), .B(N4371));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2654 (.Y(N4384), .A(N8202), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2659 (.Y(N4389), .A(N8445), .B(N8521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2660 (.Y(N6172), .A(N8213), .B(N8325));
NAND2XL hyperpropagate_3_1_A_I7423 (.Y(N8635), .A(N8354), .B(N8411));
NOR2XL hyperpropagate_3_1_A_I7424 (.Y(N4393), .A(N4384), .B(N8635));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5774 (.Y(N4396), .A(N8500), .B(N8460), .C(N4393));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5775 (.Y(N4401), .AN(N8421), .BN(N8299), .C(N4389), .D(N6172));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I10062 (.Y(N4400), .AN(N8242), .B(N133), .C(N4396), .D(N4298));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2672 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[4]), .A(N4401), .B(N4400));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2680 (.Y(N4410), .A(N8486), .B(N8247));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5778 (.Y(N6797), .AN(N164), .B(N8375));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2683 (.Y(N4413), .A(N8513), .B(N8198));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2685 (.Y(N4415), .A(N151), .B(N4410));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2686 (.Y(N4416), .A(N8315), .B(N8256));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2687 (.Y(N6799), .A(N8474), .B(N8346));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2689 (.Y(N4419), .A(N8397), .B(N8547));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5514 (.Y(N8575), .A(N8284));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2691 (.Y(N4421), .A(N8575), .B(N4413));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2692 (.Y(N4422), .A(N4419), .B(N6799));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2695 (.Y(N4425), .A(N4415), .B(N4422));
NAND3XL hyperpropagate_4_1_A_I7425 (.Y(N8644), .A(N8521), .B(N6739), .C(N4421));
NOR2XL hyperpropagate_4_1_A_I7426 (.Y(N4429), .A(N6797), .B(N8644));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I7175 (.Y(N4428), .AN(N8223), .BN(N8439), .C(N4416), .D(N4425));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2700 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[5]), .A(N4429), .B(N4428));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2705 (.Y(N4436), .A(N8168), .B(N8486));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2707 (.Y(N4438), .A(N8202), .B(N8505));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2711 (.Y(N4442), .A(N8439), .B(N8238));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2712 (.Y(N4443), .A(N8427), .B(N8372));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5788 (.Y(N4444), .AN(N8248), .B(N8379));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2714 (.Y(N6344), .A(N8186), .B(N8417));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2715 (.Y(N4446), .A(N8449), .B(N8459));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2717 (.Y(N4448), .A(N8332), .B(N8525));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2718 (.Y(N4449), .A(N6739), .B(N8213));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2720 (.Y(N4451), .A(N4438), .B(N4444));
NAND2XL hyperpropagate_3_1_A_I7427 (.Y(N8650), .A(N8366), .B(N8543));
NOR2XL hyperpropagate_3_1_A_I7428 (.Y(N4452), .A(N4449), .B(N8650));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I7177 (.Y(N4454), .AN(N146), .BN(N4436), .C(N8284), .D(N8260));
NAND2XL hyperpropagate_3_1_A_I7429 (.Y(N8657), .A(N8354), .B(N8299));
NOR2XL hyperpropagate_3_1_A_I7430 (.Y(N4455), .A(N4443), .B(N8657));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2725 (.Y(N4456), .A(N4448), .B(N6344));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2728 (.Y(N4459), .A(N4455), .B(N4456));
NAND2XL hyperpropagate_3_1_A_I7431 (.Y(N8664), .A(N4451), .B(N4452));
NOR2XL hyperpropagate_3_1_A_I7432 (.Y(N4460), .A(N4454), .B(N8664));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5797 (.Y(N4462), .A(N4446), .B(N4442), .C(N4459));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2732 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[6]), .A(N4460), .B(N4462));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2739 (.Y(N4471), .A(N133), .B(N6669));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2741 (.Y(N6356), .A(N8198), .B(N8250));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2743 (.Y(N4475), .A(N8346), .B(N8521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2744 (.Y(N6801), .A(N8383), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2745 (.Y(N4477), .A(N6739), .B(N6755));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I5799 (.Y(N8579), .A(N8482), .B(N8219));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2747 (.Y(N6805), .A(N8390), .B(N8397));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2748 (.Y(N4480), .A(N6769), .B(N8325));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2749 (.Y(N4481), .A(N6753), .B(N8546));
NAND2XL hyperpropagate_3_1_A_I7433 (.Y(N8671), .A(N8182), .B(N8264));
NOR2XL hyperpropagate_3_1_A_I7434 (.Y(N4484), .A(N6805), .B(N8671));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2753 (.Y(N4485), .A(N4480), .B(N8579));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2754 (.Y(N4486), .A(N4481), .B(N4477));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2756 (.Y(N4488), .A(N4471), .B(N4484));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5802 (.Y(N4491), .A(N4490), .B(N8575), .C(N6801));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5803 (.Y(N4493), .A(N6356), .B(N4475), .C(N4488));
NAND2XL hyperpropagate_3_1_A_I7435 (.Y(N8678), .A(N4485), .B(N4486));
NOR2XL hyperpropagate_3_1_A_I7436 (.Y(N4494), .A(N4491), .B(N8678));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2763 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[7]), .A(N4493), .B(N4494));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2768 (.Y(N4500), .A(N8411), .B(N8242));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2769 (.Y(N6807), .A(N8174), .B(N8308));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2771 (.Y(N4503), .A(N6721), .B(N6807));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2773 (.Y(N6142), .A(N8372), .B(N8379));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2774 (.Y(N5900), .A(N8182), .B(N8394));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2775 (.Y(N4507), .A(N8227), .B(N8449));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2778 (.Y(N4897), .A(N6777), .B(N8481));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2779 (.Y(N4511), .A(N8397), .B(N8260));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2782 (.Y(N4514), .A(N8575), .B(N4500));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2783 (.Y(N4515), .A(N4438), .B(N4897));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2784 (.Y(N4516), .A(N4511), .B(N4507));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2785 (.Y(N4517), .A(N6142), .B(N4481));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5806 (.Y(N4521), .A(N8460), .B(N6743), .C(N4517));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2790 (.Y(N4522), .A(N4514), .B(N4503));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6432 (.Y(N4528), .AN(N8439), .BN(N8426), .C(N5900), .D(N4475));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5808 (.Y(N4527), .AN(N4515), .BN(N4516), .C(N4522), .D(N4521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2797 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[8]), .A(N4528), .B(N4527));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2802 (.Y(N4534), .A(N8455), .B(N8198));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2803 (.Y(N4535), .A(N8426), .B(N8249));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2804 (.Y(N6531), .A(N8379), .B(N8182));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2805 (.Y(N4537), .A(N8394), .B(N8227));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2806 (.Y(N4538), .A(N8176), .B(N8288));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2807 (.Y(N4539), .A(N8402), .B(N8362));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2809 (.Y(N4541), .A(N8264), .B(N8311));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2810 (.Y(N4542), .A(N8445), .B(N8332));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2811 (.Y(N4948), .A(N6733), .B(N6739));
NAND2XL hyperpropagate_3_1_A_I7437 (.Y(N8685), .A(N8319), .B(N8350));
NOR2XL hyperpropagate_3_1_A_I7438 (.Y(N4550), .A(N4538), .B(N8685));
NAND2XL hyperpropagate_3_1_A_I7439 (.Y(N8692), .A(N8417), .B(N8210));
NOR2XL hyperpropagate_3_1_A_I7440 (.Y(N4554), .A(N4541), .B(N8692));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2816 (.Y(N4548), .A(N6791), .B(N4948));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2817 (.Y(N4549), .A(N4537), .B(N4539));
NAND2XL hyperpropagate_3_1_A_I7441 (.Y(N8699), .A(N8481), .B(N8462));
NOR2XL hyperpropagate_3_1_A_I7442 (.Y(N4552), .A(N4542), .B(N8699));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2821 (.Y(N4553), .A(N4534), .B(N6531));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2823 (.Y(N4555), .A(N4554), .B(N4535));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2824 (.Y(N4556), .A(N4548), .B(N4549));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2825 (.Y(N4560), .A(N4552), .B(N4553));
NAND3XL hyperpropagate_3_1_A_I10064 (.Y(N8706), .A(N8371), .B(N8505), .C(N4550));
NOR2XL hyperpropagate_3_1_A_I7444 (.Y(N4562), .A(N4556), .B(N8706));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2829 (.Y(N4561), .A(N4560), .B(N4555));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2831 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[9]), .A(N4562), .B(N4561));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2838 (.Y(N4591), .A(N6689), .B(N153));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2841 (.Y(N4574), .A(N8234), .B(N8513));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2842 (.Y(N4575), .A(N8372), .B(N8394));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2843 (.Y(N4576), .A(N8402), .B(N8185));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2848 (.Y(N6316), .A(N6727), .B(N8281));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2852 (.Y(N4585), .A(N6316), .B(N6799));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2853 (.Y(N4586), .A(N6797));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5822 (.Y(N4587), .AN(N4574), .B(N6769), .C(N4586));
NAND2XL hyperpropagate_3_1_A_I7445 (.Y(N8713), .A(N8417), .B(N8315));
NOR2XL hyperpropagate_3_1_A_I7446 (.Y(N4588), .A(N8579), .B(N8713));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2856 (.Y(N4589), .A(N4575), .B(N4576));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2857 (.Y(N4590), .A(N4347), .B(N5779));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2861 (.Y(N4594), .A(N4589), .B(N4590));
NAND3XL hyperpropagate_4_1_A_I7447 (.Y(N8722), .A(N4591), .B(N8332), .C(N8429));
NOR2XL hyperpropagate_4_1_A_I7448 (.Y(N4597), .A(N4594), .B(N8722));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I7196 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[10]), .AN(N4587), .B(N4588), .C(N4597), .D(N4585));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2869 (.Y(N4603), .A(N8223), .B(N8174));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5828 (.Y(N4607), .A(N8467), .B(N8439), .C(N8247));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2874 (.Y(N4608), .A(N8238), .B(N8512));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2875 (.Y(N4609), .A(N8198), .B(N8182));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2876 (.Y(N4610), .A(N8401), .B(N8210));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2880 (.Y(N4614), .A(N8383), .B(N6777));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2881 (.Y(N6809), .A(N8481), .B(N8390));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2882 (.Y(N6811), .A(N8413), .B(N6769));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2883 (.Y(N4621), .A(N8259), .B(N8546));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2884 (.Y(N4618), .A(N8470), .B(N8284));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5585 (.Y(N4625), .A(N4614), .B(N6811), .C(N6809));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I10065 (.Y(N4627), .AN(N6743), .B(N8428), .C(N4608), .D(N4609));
NAND2XL hyperpropagate_3_1_A_I7449 (.Y(N8728), .A(N8315), .B(N8366));
NOR2XL hyperpropagate_3_1_A_I7450 (.Y(N4628), .A(N4610), .B(N8728));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5835 (.Y(N4634), .A(N4603), .B(N4618), .C(N4448));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6450 (.Y(N4631), .A(N6697), .B(N6705), .C(N4621), .D(N4607));
NAND2XL hyperpropagate_3_1_A_I7451 (.Y(N8735), .A(N4628), .B(N4625));
NOR2XL hyperpropagate_3_1_A_I7452 (.Y(N4635), .A(N4634), .B(N8735));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I10067 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[11]), .A(N4631), .B(N4627), .C(N4635));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2909 (.Y(N4643), .A(N8202), .B(N8486));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2911 (.Y(N4645), .A(N8478), .B(N8407));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2913 (.Y(N4647), .A(N8421), .B(N8238));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5845 (.Y(N4652), .A(N8354), .B(N8174), .C(N8332));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2919 (.Y(N6813), .A(N8509), .B(N6739));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2920 (.Y(N4654), .A(N6755), .B(N8281));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I2921 (.Y(N6815), .A(N8324), .B(N6753));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2922 (.Y(N4656), .A(N8546));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5846 (.Y(N4659), .A(N4645), .B(N4643), .C(N6815));
NAND2XL hyperpropagate_3_1_A_I7453 (.Y(N8742), .A(N8535), .B(N8256));
NOR2XL hyperpropagate_3_1_A_I7454 (.Y(N4661), .A(N6344), .B(N8742));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5850 (.Y(N4669), .A(N4652), .B(N6797), .C(N6813));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2932 (.Y(N4667), .A(N4659), .B(N4661));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I10068 (.Y(N4668), .A(N4656), .B(N4647), .C(N4654), .D(N4667));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2936 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[12]), .A(N4669), .B(N4668));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2942 (.Y(N4677), .A(N8247), .B(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2943 (.Y(N4678), .A(N8411), .B(N8174));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2947 (.Y(N4682), .A(N128), .B(N4677));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5853 (.Y(N4684), .A(N8467), .B(N8486), .C(N8421));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2950 (.Y(N4685), .A(N8455), .B(N8496));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2951 (.Y(N4686), .A(N8372), .B(N8182));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2953 (.Y(N4688), .A(N8366), .B(N8474));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2954 (.Y(N4689), .A(N8346));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5855 (.Y(N4692), .A(N8288), .B(N8332), .C(N8264));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2959 (.Y(N6817), .A(N8218), .B(N8390));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2961 (.Y(N4696), .A(N8324));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2962 (.Y(N4697), .A(N4696), .B(N4688));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2963 (.Y(N4702), .A(N4678), .B(N6817));
NAND2XL hyperpropagate_3_1_A_I7455 (.Y(N8749), .A(N8397), .B(N8213));
NOR2XL hyperpropagate_3_1_A_I7456 (.Y(N4699), .A(N6813), .B(N8749));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I7204 (.Y(N4708), .A(N8202), .B(N8299), .C(N4697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2969 (.Y(N4704), .A(N4682), .B(N4699));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5859 (.Y(N4706), .A(N4684), .B(N4685), .C(N4689));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2972 (.Y(N4707), .A(N4692), .B(N4704));
NAND3XL hyperpropagate_4_1_A_I10095 (.Y(N11621), .A(N4702), .B(N4686), .C(N4706));
NOR2XL hyperpropagate_4_1_A_I10096 (.Y(N4710), .A(N4708), .B(N11621));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2976 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[13]), .A(N4710), .B(N4707));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2983 (.Y(N4718), .A(N8247), .B(N8319));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2984 (.Y(N4719), .A(N8354), .B(N8308));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5866 (.Y(N4733), .AN(N160), .B(N8168), .C(N8539));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2988 (.Y(N4723), .A(N8512), .B(N8496));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2989 (.Y(N4724), .A(N8551), .B(N8427));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2991 (.Y(N4737), .A(N8521), .B(N8383));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2992 (.Y(N5610), .A(N6727), .B(N8481));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2996 (.Y(N4731), .A(N4298), .B(N6811));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2997 (.Y(N4732), .A(N4718), .B(N4719));
NAND2XL hyperpropagate_3_1_A_I7457 (.Y(N8756), .A(N8227), .B(N8210));
NOR2XL hyperpropagate_3_1_A_I7458 (.Y(N4735), .A(N4723), .B(N8756));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3001 (.Y(N4736), .A(N5610), .B(N4724));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5869 (.Y(N4740), .A(N8299), .B(N8233), .C(N4735));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3006 (.Y(N4741), .A(N4731), .B(N4736));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I7208 (.Y(N4743), .A(N4733), .B(N6805), .C(N4741));
NAND2XL hyperpropagate_3_1_A_I7459 (.Y(N8763), .A(N4737), .B(N4732));
NOR2XL hyperpropagate_3_1_A_I7460 (.Y(N4744), .A(N4740), .B(N8763));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3010 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[14]), .A(N4743), .B(N4744));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3018 (.Y(N5300), .A(N8350), .B(N8206));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3019 (.Y(N4755), .A(N8238), .B(N8500));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5874 (.Y(N8594), .A(N8512), .B(N8277));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5534 (.Y(N8595), .A(N8594));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3022 (.Y(N4769), .A(N8264), .B(N8315));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I6473 (.Y(N8598), .A(N8462), .B(N6753));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3026 (.Y(N4762), .A(N8546), .B(N8515));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3027 (.Y(N4767), .A(N6697), .B(N5300));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3029 (.Y(N4765), .A(N8598), .B(N6316));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I7212 (.Y(N4772), .A(N8482), .B(N6769), .C(N4767));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6476 (.Y(N4774), .AN(N8250), .BN(N8227), .C(N4762), .D(N4769));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I7213 (.Y(N4771), .AN(N4755), .B(N8594), .C(N4765));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3037 (.Y(N4773), .A(N4772), .B(N4771));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3039 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[15]), .A(N4774), .B(N4773));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I6479 (.Y(N4778), .AN(N144), .B(N8371));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3048 (.Y(N4784), .A(N8350), .B(N8407));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3053 (.Y(N4789), .A(N8459), .B(N8366));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3054 (.Y(N4790), .A(N8255), .B(N8474));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3058 (.Y(N4794), .A(N8525), .B(N8509));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3059 (.Y(N4795), .A(N6727), .B(N8213));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3061 (.Y(N4805), .A(N4290), .B(N4444));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I7214 (.Y(N4799), .AN(N8500), .BN(N8277), .C(N4794), .D(N4795));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I7215 (.Y(N4801), .AN(N8486), .BN(N8435), .C(N4789), .D(N4784));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3066 (.Y(N4802), .A(N4724), .B(N4790));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5890 (.Y(N4804), .A(N149), .B(N4778), .C(N4347));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I10070 (.Y(N4809), .A(N8449), .B(N8332), .C(N8288), .D(N4805));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3071 (.Y(N4807), .A(N4802), .B(N4799));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3074 (.Y(N4810), .A(N4809), .B(N4807));
NAND3X1 inst_cellmath__195__80__2WWMM_2WWMM_I10072 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[16]), .A(N4804), .B(N4801), .C(N4810));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3084 (.Y(N4821), .A(N8130), .B(N6711));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3085 (.Y(N4822), .A(N8354), .B(N8528));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3087 (.Y(N4824), .A(N8250), .B(N8176));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3088 (.Y(N4825), .A(N8449), .B(N8366));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3089 (.Y(N4826), .A(N8474), .B(N8311));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3090 (.Y(N4827), .A(N8445), .B(N4821));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I5897 (.Y(N4829), .AN(N4824), .B(N8332));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3093 (.Y(N4839), .A(N8521), .B(N6777));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3094 (.Y(N4831), .A(N6755), .B(N8390));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3095 (.Y(N4832), .A(N8189), .B(N8413));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3098 (.Y(N4835), .A(N4831), .B(N4827));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I7320 (.Y(N4842), .AN(N4825), .BN(N4826), .C(N8299), .D(N8512));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I7220 (.Y(N4847), .AN(N8259), .B(N4822), .C(N4829), .D(N4832));
NAND2XL hyperpropagate_3_1_A_I7461 (.Y(N8770), .A(N4839), .B(N4835));
NOR2XL hyperpropagate_3_1_A_I7462 (.Y(N4846), .A(N4842), .B(N8770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3111 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[17]), .A(N4847), .B(N4846));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3122 (.Y(N4860), .A(N6719), .B(N6695));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3123 (.Y(N6278), .A(N8455), .B(N8512));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6497 (.Y(N4865), .A(N8444), .B(N8362), .C(N8250), .D(N4860));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3128 (.Y(N4866), .A(N8332), .B(N6739));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5908 (.Y(N4875), .A(N6809), .B(N6278), .C(N4865));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6499 (.Y(N4876), .A(N6795), .B(N4511), .C(N6799), .D(N4866));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3139 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[18]), .A(N4875), .B(N4876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3148 (.Y(N4886), .A(N8505), .B(N8339));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3149 (.Y(N4887), .A(N8250), .B(N6743));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3154 (.Y(N6563), .A(N8413), .B(N8259));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3155 (.Y(N4893), .A(N8324), .B(N8284));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5912 (.Y(N4901), .AN(N6805), .B(N8430), .C(N6739));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5914 (.Y(N4900), .A(N4886), .B(N4826), .C(N4887));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I5916 (.Y(N4902), .A(N4893), .B(N4897), .C(N6563), .D(N4901));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3165 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[19]), .A(N4900), .B(N4902));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3176 (.Y(N6823), .A(N8444), .B(N8430));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3177 (.Y(N4915), .A(N6733), .B(N6727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3179 (.Y(N4917), .A(N8397), .B(N8189));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3181 (.Y(N4919), .A(N8213), .B(N8462));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3184 (.Y(N4922), .A(N6811), .B(N6817));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6500 (.Y(N4924), .AN(N8478), .BN(N8176), .C(N4917), .D(N4919));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I5922 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[20]), .AN(N4915), .BN(N6823), .C(N4922), .D(N4924));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3199 (.Y(N4937), .A(N8346), .B(N8383));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3202 (.Y(N4940), .A(N8218), .B(N8189));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I6501 (.Y(N8601), .A(N8212), .B(N8259));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5542 (.Y(N8603), .A(N8601));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I5541 (.Y(N8602), .A(N8601));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3205 (.Y(N4943), .A(N8336), .B(N8284));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3207 (.Y(N4945), .A(N4940), .B(N8603));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3208 (.Y(N4946), .A(N6815), .B(N4943));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I7223 (.Y(N4953), .AN(N6743), .BN(N8311), .C(N6789), .D(N4948));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3212 (.Y(N4950), .A(N4945), .B(N4946));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5926 (.Y(N4952), .A(N4937), .B(N4824), .C(N4950));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3216 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[21]), .A(N4953), .B(N4952));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3241 (.Y(N4979), .A(N8206), .B(N8427));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3242 (.Y(N4980), .A(N8379), .B(N8227));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3246 (.Y(N4984), .A(N8311), .B(N8346));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3253 (.Y(N4991), .A(N8470));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3254 (.Y(N4992), .A(N4991), .B(N4980));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6506 (.Y(N4995), .A(N8481), .B(N8546), .C(N8255), .D(N8366));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3260 (.Y(N4998), .A(N4839), .B(N4992));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I7463 (.Y(N8779), .A(N8386), .B(N8299), .C(N8129));
NAND3XL hyperpropagate_4_1_A_I7465 (.Y(N8787), .A(N8445), .B(N8247), .C(N8411));
NOR4X1 hyperpropagate_4_1_A_I10073 (.Y(N5002), .A(N4979), .B(N6787), .C(N4993), .D(N8787));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I10074 (.Y(N5005), .AN(N5002), .B(N8779), .C(N4995));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I5936 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[23]), .AN(N4984), .BN(N4998), .C(N8332), .D(N5005));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3276 (.Y(N5014), .A(N8467), .B(N8294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5938 (.Y(N8605), .A(N8505), .B(N8435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3279 (.Y(N5017), .A(N8407), .B(N8455));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3281 (.Y(N5019), .A(N6715), .B(N5014));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3282 (.Y(N5020), .A(N8372), .B(N8249));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3283 (.Y(N6139), .A(N8487), .B(N8394));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3287 (.Y(N5025), .A(N8189), .B(N8324));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5940 (.Y(N5031), .AN(N5025), .B(N8543), .C(N5019), .D(N8430));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6507 (.Y(N5038), .AN(N6139), .BN(N4603), .C(N8255), .D(N8362));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6508 (.Y(N5036), .A(N5017), .B(N8605), .C(N8575), .D(N5020));
NAND2XL hyperpropagate_3_1_A_I7467 (.Y(N8793), .A(N8521), .B(N6733));
NOR2XL hyperpropagate_3_1_A_I7468 (.Y(N5035), .A(N5031), .B(N8793));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5946 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[24]), .AN(N5038), .B(N5036), .C(N5035));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3316 (.Y(N5055), .A(N8417), .B(N8535));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3317 (.Y(N5056), .A(N8474), .B(N8444));
NAND2XL hyperpropagate_3_1_A_I7469 (.Y(N8800), .A(N8294), .B(N8486));
NOR2XL hyperpropagate_3_1_A_I7470 (.Y(N5061), .A(N4348), .B(N8800));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I5950 (.Y(N5063), .A(N8319), .B(N8462), .C(N8339), .D(N5061));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6510 (.Y(N5065), .AN(N8372), .BN(N8401), .C(N6679), .D(N112));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5952 (.Y(N5067), .AN(N8218), .BN(N8259), .C(N5055), .D(N5056));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3330 (.Y(N5069), .A(N5065), .B(N5067));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5955 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[25]), .AN(N5063), .B(N8281), .C(N5069), .D(N8521));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3339 (.Y(N5078), .A(N8486), .B(N8354));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3342 (.Y(N5081), .A(N8198), .B(N8551));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5957 (.Y(N8607), .A(N8336), .B(N8515));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5958 (.Y(N5090), .AN(N5078), .B(N8210), .C(N8366));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6729 (.Y(N5099), .AN(N6739), .BN(N8325), .C(N8607), .D(N6801));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3357 (.Y(N5096), .A(N4723), .B(N4575));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5963 (.Y(N5098), .AN(N8288), .BN(N8185), .C(N4790), .D(N5081));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I5964 (.Y(N5102), .AN(N5090), .B(N8304), .C(N5098), .D(N8407));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I5965 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[26]), .AN(N5102), .B(N5096), .C(N5099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3370 (.Y(N5110), .A(N8539), .B(N8319));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3371 (.Y(N5126), .A(N8308), .B(N8350));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3376 (.Y(N5116), .A(N8394), .B(N8401));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3377 (.Y(N5128), .A(N8417), .B(N8264));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I5967 (.Y(N8609), .A(N8547), .B(N8470));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5968 (.Y(N5127), .A(N122), .B(N6695), .C(N5126));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5969 (.Y(N5129), .A(N8567), .B(N5128), .C(N8609));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6512 (.Y(N5131), .AN(N5110), .BN(N4940), .C(N8508), .D(N8482));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3392 (.Y(N5135), .A(N5116), .B(N4789));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3394 (.Y(N5134), .A(N5127), .B(N5129));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3396 (.Y(N5136), .A(N5135), .B(N4737));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I7224 (.Y(N5140), .AN(N8198), .BN(N8427), .C(N5020), .D(N5131));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3399 (.Y(N5139), .A(N5134), .B(N5136));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3401 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[27]), .A(N5140), .B(N5139));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3408 (.Y(N5148), .A(N8371), .B(N8294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3415 (.Y(N5155), .A(N8535), .B(N8315));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3416 (.Y(N5156), .A(N8459), .B(N8255));
AND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5976 (.Y(N5172), .A(N8304), .B(N8332), .C(N8247));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3419 (.Y(N5163), .A(N8383), .B(N8281));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3421 (.Y(N5161), .A(N8413), .B(N6753));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5977 (.Y(N5164), .A(N155), .B(N5163), .C(N5148));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6516 (.Y(N5167), .AN(N8198), .BN(N8185), .C(N6817), .D(N5161));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3428 (.Y(N5168), .A(N4723), .B(N5156));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5979 (.Y(N5170), .A(N4292), .B(N5155), .C(N5164));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6517 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[28]), .A(N5172), .B(N5168), .C(N5167), .D(N5170));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3443 (.Y(N5184), .A(N8386), .B(N8247));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3444 (.Y(N5185), .A(N8299), .B(N8407));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3449 (.Y(N5190), .A(N8315), .B(N8346));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3450 (.Y(N5198), .A(N8445), .B(N8482));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5986 (.Y(N5205), .AN(N6769), .BN(N6753), .C(N5184), .D(N5198));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I5987 (.Y(N5201), .A(N8575), .B(N6791), .C(N5190));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5988 (.Y(N5203), .AN(N8233), .BN(N8500), .C(N4351), .D(N5128));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3463 (.Y(N5204), .A(N5185), .B(N8595));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6518 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[29]), .A(N5203), .B(N5201), .C(N5205), .D(N5204));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3476 (.Y(N5218), .A(N8223), .B(N8308));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3481 (.Y(N5223), .A(N8459), .B(N8543));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3482 (.Y(N5224), .A(N6743), .B(N8525));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3483 (.Y(N5225), .A(N6739), .B(N6727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3484 (.Y(N5226), .A(N6755), .B(N6769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3487 (.Y(N5229), .A(N4696), .B(N5224));
NAND2XL hyperpropagate_3_1_A_I7471 (.Y(N8807), .A(N8487), .B(N8288));
NOR2XL hyperpropagate_3_1_A_I7472 (.Y(N5230), .A(N5226), .B(N8807));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3494 (.Y(N5236), .A(N4586), .B(N5229));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6520 (.Y(N5238), .AN(N8401), .BN(N8417), .C(N5218), .D(N8602));
NAND3XL hyperpropagate_4_1_A_I7473 (.Y(N8816), .A(N8478), .B(N8421), .C(N5225));
NOR2XL hyperpropagate_4_1_A_I7474 (.Y(N5240), .A(N5223), .B(N8816));
NAND3XL hyperpropagate_4_1_A_I7475 (.Y(N8824), .A(N8539), .B(N8247), .C(N5230));
NOR2XL hyperpropagate_4_1_A_I7476 (.Y(N5243), .A(N5236), .B(N8824));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I5999 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[30]), .A(N5238), .B(N5243), .C(N5240));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3511 (.Y(N6833), .A(N8426), .B(N8379));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3513 (.Y(N5264), .A(N8449), .B(N8210));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3518 (.Y(N5260), .A(N8332), .B(N6727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3519 (.Y(N5261), .A(N8390), .B(N8189));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3521 (.Y(N5263), .A(N4621), .B(N5261));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6001 (.Y(N5265), .AN(N4538), .B(N8486), .C(N5264), .D(N8371));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6002 (.Y(N5267), .A(N8354), .B(N8500), .C(N5263));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3527 (.Y(N5273), .A(N5056), .B(N6787));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3528 (.Y(N5270), .A(N8595), .B(N5265));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6733 (.Y(N5272), .AN(N8366), .BN(N6743), .C(N6833), .D(N5267));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6524 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[31]), .A(N5260), .B(N5273), .C(N5272), .D(N5270));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3542 (.Y(N5927), .A(N8411), .B(N8339));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3543 (.Y(N5285), .A(N8242), .B(N8174));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I6007 (.Y(N5287), .AN(N4778), .B(N8299));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3550 (.Y(N5302), .A(N8185), .B(N8535));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3552 (.Y(N5294), .A(N138), .B(N5285));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3553 (.Y(N5306), .A(N8255), .B(N8310));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6525 (.Y(N5298), .A(N8470), .B(N8324), .C(N8383), .D(N8464));
NAND3XL hyperpropagate_4_1_A_I7477 (.Y(N8832), .A(N8288), .B(N8551), .C(N5927));
NOR2XL hyperpropagate_4_1_A_I7478 (.Y(N5308), .A(N5302), .B(N8832));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6526 (.Y(N5304), .A(N8421), .B(N8455), .C(N8198), .D(N8277));
NAND2XL hyperpropagate_3_1_A_I7479 (.Y(N8838), .A(N5306), .B(N5304));
NOR4X1 hyperpropagate_3_1_A_I10075 (.Y(N5311), .A(N5300), .B(N5298), .C(N5287), .D(N8838));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6017 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[32]), .A(N5294), .B(N5308), .C(N5311));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3579 (.Y(N5321), .A(N8304), .B(N8206));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3582 (.Y(N5324), .A(N8315), .B(N6743));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3585 (.Y(N5335), .A(N8482), .B(N8188));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6734 (.Y(N5330), .A(N6769), .B(N8260), .C(N8336), .D(N8464));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3589 (.Y(N5331), .A(N8605), .B(N4654));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6022 (.Y(N5339), .AN(N8223), .BN(N8528), .C(N5321), .D(N5324));
NAND3XL hyperpropagate_4_1_A_I7481 (.Y(N8847), .A(N8247), .B(N8129), .C(N5330));
NOR2XL hyperpropagate_4_1_A_I7482 (.Y(N5340), .A(N6799), .B(N8847));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6528 (.Y(N5342), .AN(N5335), .BN(N5331), .C(N4755), .D(N5116));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6025 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[33]), .A(N5339), .B(N5340), .C(N5342));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3608 (.Y(N5350), .A(N8129), .B(N8294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3611 (.Y(N5353), .A(N8242), .B(N8478));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3613 (.Y(N5355), .A(N8238), .B(N8496));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3616 (.Y(N5358), .A(N123), .B(N5350));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3621 (.Y(N5363), .A(N8255), .B(N8430));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3624 (.Y(N5366), .A(N5161), .B(N5355));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6028 (.Y(N5368), .AN(N8539), .BN(N8505), .C(N4778), .D(N5353));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3627 (.Y(N5369), .A(N4980), .B(N5321));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3628 (.Y(N5370), .A(N5366), .B(N5358));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3629 (.Y(N5371), .A(N5369), .B(N5368));
NAND3XL hyperpropagate_4_1_A_I7483 (.Y(N8855), .A(N8459), .B(N8319), .C(N8435));
NOR2XL hyperpropagate_4_1_A_I7484 (.Y(N5376), .A(N5363), .B(N8855));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3632 (.Y(N5374), .A(N5370), .B(N5371));
NAND3XL hyperpropagate_4_1_A_I7485 (.Y(N8863), .A(N8521), .B(N6727), .C(N5376));
NOR2XL hyperpropagate_4_1_A_I7486 (.Y(N5375), .A(N4993), .B(N8863));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3635 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[34]), .A(N5374), .B(N5375));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3643 (.Y(N5385), .A(N8435), .B(N8350));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6531 (.Y(N5394), .AN(N8310), .BN(N8429), .C(N163), .D(N5350));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I6035 (.Y(N5396), .AN(N5385), .B(N8332));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3657 (.Y(N5399), .A(N8464), .B(N8515));
NAND2XL hyperpropagate_3_1_A_I7487 (.Y(N8869), .A(N8218), .B(N8413));
NOR2XL hyperpropagate_3_1_A_I7488 (.Y(N5402), .A(N5399), .B(N8869));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3664 (.Y(N5406), .A(N4688), .B(N4610));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6041 (.Y(N5410), .AN(N5406), .B(N5163), .C(N4769), .D(N5355));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6042 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[35]), .AN(N5396), .B(N5402), .C(N5410), .D(N5394));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3677 (.Y(N5420), .A(N8277), .B(N8426));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3680 (.Y(N5423), .A(N8535));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3684 (.Y(N5427), .A(N8346), .B(N8444));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3686 (.Y(N5429), .A(N8188), .B(N8212));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3687 (.Y(N6354), .A(N8325), .B(N8547));
NAND2XL hyperpropagate_3_1_A_I7489 (.Y(N8876), .A(N8478), .B(N8238));
NOR2XL hyperpropagate_3_1_A_I7490 (.Y(N5439), .A(N5427), .B(N8876));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6533 (.Y(N5435), .A(N5429), .B(N6705), .C(N5423), .D(N6795));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6048 (.Y(N5438), .AN(N6354), .B(N6727), .C(N5420), .D(N8218));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6050 (.Y(N5442), .AN(N6139), .B(N8449), .C(N4586), .D(N8176));
NAND3XL hyperpropagate_4_1_A_I7491 (.Y(N8885), .A(N8460), .B(N8411), .C(N8294));
NOR2XL hyperpropagate_4_1_A_I7492 (.Y(N5447), .A(N5438), .B(N8885));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6537 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[36]), .AN(N5442), .B(N5439), .C(N5447), .D(N5435));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3710 (.Y(N5454), .A(N8202), .B(N8168));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3717 (.Y(N5461), .A(N8206), .B(N8375));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3721 (.Y(N5465), .A(N8449), .B(N8264));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3722 (.Y(N5466), .A(N8430));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6538 (.Y(N5467), .AN(N8182), .B(N6711), .C(N5466), .D(N5454));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3727 (.Y(N6212), .A(N6733), .B(N8508));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3728 (.Y(N6835), .A(N6777), .B(N6755));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3730 (.Y(N5474), .A(N124), .B(N6835));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6057 (.Y(N5482), .AN(N8319), .BN(N8242), .C(N5465), .D(N5461));
NAND3XL hyperpropagate_4_1_A_I7493 (.Y(N8893), .A(N8277), .B(N8487), .C(N5467));
NOR2XL hyperpropagate_4_1_A_I7494 (.Y(N5481), .A(N4539), .B(N8893));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6060 (.Y(N5486), .AN(N6212), .BN(N5126), .C(N5474), .D(N5482));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6061 (.Y(N5485), .A(N8386), .B(N8332), .C(N8223), .D(N5481));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3743 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[37]), .A(N5486), .B(N5485));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3753 (.Y(N5497), .A(N8242), .B(N8277));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3754 (.Y(N5498), .A(N8379), .B(N8178));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3760 (.Y(N5508), .A(N6755), .B(N8218));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3761 (.Y(N5505), .A(N8413), .B(N8464));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3763 (.Y(N5507), .A(N4991), .B(N5505));
NAND3XL hyperpropagate_4_1_A_I7495 (.Y(N8901), .A(N8310), .B(N5508), .C(N5507));
NOR2XL hyperpropagate_4_1_A_I7496 (.Y(N5512), .A(N5078), .B(N8901));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6066 (.Y(N5517), .AN(N8255), .BN(N8449), .C(N5498), .D(N5497));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3774 (.Y(N5518), .A(N5517), .B(N5260));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6916 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[38]), .AN(N5518), .B(N8288), .C(N5512), .D(N8401));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3795 (.Y(N5539), .A(N6753), .B(N8284));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6542 (.Y(N5545), .AN(N6733), .BN(N8218), .C(N5539), .D(N4832));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6741 (.Y(N5544), .AN(N8277), .BN(N8178), .C(N5466), .D(N5427));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6917 (.Y(N5547), .A(N8401), .B(N8332), .C(N6743), .D(N8455));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6077 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[39]), .A(N8247), .B(N5545), .C(N5544), .D(N5547));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3815 (.Y(N5560), .A(N8310), .B(N8444));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3817 (.Y(N5562), .A(N6777), .B(N6727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3821 (.Y(N5566), .A(N8464), .B(N8547));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6079 (.Y(N5570), .AN(N5566), .B(N8535), .C(N6743));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3826 (.Y(N5575), .A(N6791), .B(N5560));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3827 (.Y(N5572), .A(N6172), .B(N5562));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6080 (.Y(N5574), .AN(N6811), .B(N8277), .C(N8339));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3831 (.Y(N5576), .A(N5575), .B(N5335));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6081 (.Y(N5579), .AN(N8575), .B(N8429), .C(N5572), .D(N8508));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3835 (.Y(N5583), .A(N5579), .B(N5576));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6547 (.Y(N5582), .AN(N8178), .BN(N8401), .C(N5574), .D(N5570));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3839 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[40]), .A(N5583), .B(N5582));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6548 (.Y(N5593), .A(N8401), .B(N8176), .C(N8129), .D(N8249));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3849 (.Y(N5594), .A(N8535), .B(N8445));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3850 (.Y(N5595), .A(N8429), .B(N6733));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3851 (.Y(N5596), .A(N8508), .B(N6777));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3859 (.Y(N5604), .A(N5566), .B(N6791));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3863 (.Y(N5608), .A(N4940));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3864 (.Y(N5609), .A(N5608), .B(N5604));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6086 (.Y(N5614), .A(N5610), .B(N5594), .C(N8602));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6549 (.Y(N5613), .A(N5595), .B(N6811), .C(N5596), .D(N5609));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6090 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[41]), .AN(N5593), .B(N5614), .C(N5613));
NAND2XL hyperpropagate_3_1_A_I7497 (.Y(N8907), .A(N8407), .B(N8249));
NOR2XL hyperpropagate_3_1_A_I7498 (.Y(N5635), .A(N5261), .B(N8907));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3893 (.Y(N5641), .A(N5225), .B(N5508));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6093 (.Y(N5639), .AN(N6801), .B(N8178), .C(N5635), .D(N6743));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6550 (.Y(N5643), .A(N6815), .B(N4943), .C(N4984), .D(N8602));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3897 (.Y(N5642), .A(N5641), .B(N5639));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3899 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[42]), .A(N5643), .B(N5642));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3908 (.Y(N5654), .A(N8233), .B(N8277));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I3911 (.Y(N5657), .A(N6743));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3916 (.Y(N5662), .A(N4689), .B(N8605));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6099 (.Y(N5664), .AN(N5657), .B(N8543), .C(N8535), .D(N8247));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3919 (.Y(N5751), .A(N8332), .B(N8383));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3923 (.Y(N5669), .A(N8562), .B(N8602));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3925 (.Y(N5671), .A(N5608), .B(N5669));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6102 (.Y(N5675), .AN(N8474), .B(N6807), .C(N5664));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6103 (.Y(N5680), .AN(N8421), .BN(N8500), .C(N5654), .D(N5671));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6104 (.Y(N5682), .AN(N5662), .B(N8198), .C(N5675), .D(N8362));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6105 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[43]), .AN(N5682), .B(N5751), .C(N5680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3942 (.Y(N5689), .A(N8319), .B(N8354));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3947 (.Y(N5694), .A(N8210), .B(N6743));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3955 (.Y(N5702), .A(N6807), .B(N8607));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6552 (.Y(N5707), .A(N8218), .B(N8394), .C(N8397), .D(N8417));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6109 (.Y(N5708), .AN(N5694), .B(N8470), .C(N5702), .D(N8188));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6112 (.Y(N5713), .A(N6789), .B(N6801), .C(N5596), .D(N5708));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6113 (.Y(N5714), .AN(N6713), .BN(N5689), .C(N4535), .D(N5713));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6114 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[44]), .AN(N5714), .B(N8528), .C(N5707), .D(N8277));
NAND2XL hyperpropagate_3_1_A_I7499 (.Y(N8914), .A(N8543), .B(N8346));
NOR2XL hyperpropagate_3_1_A_I7500 (.Y(N5731), .A(N5466), .B(N8914));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3990 (.Y(N5738), .A(N6753), .B(N8470));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I3991 (.Y(N5741), .A(N4268), .B(N5738));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I3994 (.Y(N5742), .A(N5741), .B(N4686));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6553 (.Y(N5744), .AN(N8299), .BN(N8198), .C(N106), .D(N8130));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6119 (.Y(N5746), .AN(N8281), .BN(N8397), .C(N5505), .D(N4416));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6120 (.Y(N5748), .AN(N5742), .B(N8174), .C(N5731), .D(N8505));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6122 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[45]), .AN(N5748), .B(N5744), .C(N5751), .D(N5746));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4012 (.Y(N6457), .A(N8487), .B(N8182));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4019 (.Y(N5768), .A(N6769), .B(N8212));
NAND2XL hyperpropagate_3_1_A_I7501 (.Y(N8921), .A(N6733), .B(N6755));
NOR2XL hyperpropagate_3_1_A_I7502 (.Y(N5771), .A(N5560), .B(N8921));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4023 (.Y(N5772), .A(N5539), .B(N6457));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4024 (.Y(N5773), .A(N4326), .B(N91));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6125 (.Y(N5774), .AN(N5768), .B(N8429), .C(N5771), .D(N8525));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4028 (.Y(N5777), .A(N5774), .B(N5155));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6128 (.Y(N5781), .AN(N8595), .B(N5773), .C(N5777), .D(N5772));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6129 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[46]), .A(N6797), .B(N5779), .C(N5185), .D(N5781));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4041 (.Y(N5791), .A(N8168), .B(N8294));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4051 (.Y(N5801), .A(N8260), .B(N8470));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4053 (.Y(N5803), .A(N8575), .B(N5791));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4054 (.Y(N5804), .A(N4643), .B(N5110));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4055 (.Y(N5805), .A(N5801), .B(N4319));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4056 (.Y(N5806), .A(N5461), .B(N4296));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4058 (.Y(N5808), .A(N5803), .B(N5804));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4059 (.Y(N5809), .A(N5805), .B(N5806));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6132 (.Y(N5812), .AN(N8525), .BN(N8218), .C(N4719), .D(N5809));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6133 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[47]), .AN(N5808), .B(N8372), .C(N5812), .D(N8362));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4070 (.Y(N5821), .A(N8319), .B(N8174));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4072 (.Y(N5823), .A(N113), .B(N6719));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4075 (.Y(N6837), .A(N8362), .B(N8210));
NAND2XL hyperpropagate_3_1_A_I7503 (.Y(N8928), .A(N8264), .B(N8346));
NOR2XL hyperpropagate_3_1_A_I7504 (.Y(N5835), .A(N6837), .B(N8928));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6138 (.Y(N5838), .AN(N6769), .BN(N8547), .C(N4537), .D(N8607));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6139 (.Y(N5839), .AN(N5562), .B(N8445), .C(N5835), .D(N6739));
NAND3XL hyperpropagate_4_1_A_I7505 (.Y(N8937), .A(N6755), .B(N8413), .C(N5838));
NOR2XL hyperpropagate_4_1_A_I7506 (.Y(N5842), .A(N5821), .B(N8937));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6142 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[48]), .AN(N5839), .B(N5823), .C(N5842), .D(N8401));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4100 (.Y(N5865), .A(N8227), .B(N8417));
NAND2XL hyperpropagate_3_1_A_I7507 (.Y(N8943), .A(N8407), .B(N8551));
NOR2XL hyperpropagate_3_1_A_I7508 (.Y(N5853), .A(N5350), .B(N8943));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4110 (.Y(N5861), .A(N5596), .B(N5768));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4113 (.Y(N5864), .A(N6457), .B(N4444));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4115 (.Y(N5866), .A(N5865), .B(N5861));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6146 (.Y(N5869), .AN(N8598), .B(N8304), .C(N5864), .D(N8339));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4121 (.Y(N5872), .A(N5155), .B(N5869));
NAND3XL hyperpropagate_4_1_A_I7509 (.Y(N8952), .A(N6727), .B(N8390), .C(N5853));
NOR2XL hyperpropagate_4_1_A_I7510 (.Y(N5875), .A(N4790), .B(N8952));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6149 (.Y(N5874), .AN(N5872), .B(N6823), .C(N5866), .D(N6795));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4125 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[49]), .A(N5875), .B(N5874));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4132 (.Y(N5884), .A(N8247), .B(N8478));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4133 (.Y(N5885), .A(N8407), .B(N8439));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4134 (.Y(N5886), .A(N8500), .B(N8551));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4137 (.Y(N6314), .A(N8227), .B(N8178));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4140 (.Y(N5892), .A(N5423), .B(N6314));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6151 (.Y(N5906), .A(N5226), .B(N5399), .C(N5900));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6152 (.Y(N5903), .A(N6833), .B(N6713), .C(N5885));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6153 (.Y(N5908), .AN(N8288), .BN(N8210), .C(N5884), .D(N5886));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6554 (.Y(N5910), .A(N5903), .B(N5892), .C(N8332), .D(N5906));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6155 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[50]), .A(N5908), .B(N5306), .C(N5910));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4166 (.Y(N5919), .A(N6719), .B(N6679));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4175 (.Y(N5928), .A(N5927), .B(N5919));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4177 (.Y(N5930), .A(N8525), .B(N8482));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6555 (.Y(N5935), .A(N8505), .B(N8206), .C(N8319), .D(N8407));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6556 (.Y(N5936), .A(N8182), .B(N8379), .C(N8551), .D(N8227));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6160 (.Y(N5938), .AN(N8390), .BN(N8260), .C(N8575), .D(N5928));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6161 (.Y(N5939), .AN(N5930), .B(N8362), .C(N5935), .D(N6743));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4189 (.Y(N5942), .A(N6799), .B(N5939));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4190 (.Y(N5943), .A(N5938), .B(N5942));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6163 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[51]), .AN(N5943), .B(N8439), .C(N5936), .D(N8500));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6165 (.Y(N5963), .A(N6689), .B(N6669), .C(N4291));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4212 (.Y(N6065), .A(N8508), .B(N8281));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4213 (.Y(N5967), .A(N8397), .B(N6769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4216 (.Y(N5970), .A(N8562), .B(N5967));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4217 (.Y(N5971), .A(N6815), .B(N6065));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4220 (.Y(N5974), .A(N5970), .B(N5963));
NAND3XL hyperpropagate_4_1_A_I7511 (.Y(N8960), .A(N8474), .B(N8435), .C(N8129));
NOR2XL hyperpropagate_4_1_A_I7512 (.Y(N5975), .A(N5974), .B(N8960));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6168 (.Y(N5977), .AN(N5971), .B(N8206), .C(N5975), .D(N8372));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6169 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[52]), .AN(N5977), .B(N5865), .C(N8332));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4241 (.Y(N5996), .A(N6701), .B(N5385));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4243 (.Y(N5998), .A(N8188), .B(N8464));
NAND2XL hyperpropagate_3_1_A_I7513 (.Y(N8966), .A(N8233), .B(N8426));
NOR2XL hyperpropagate_3_1_A_I7514 (.Y(N6004), .A(N4575), .B(N8966));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6173 (.Y(N6006), .AN(N8539), .BN(N8500), .C(N5017), .D(N6314));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6174 (.Y(N6010), .AN(N6004), .B(N8609), .C(N5998), .D(N6837));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4256 (.Y(N6011), .A(N6010), .B(N5996));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6176 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[53]), .AN(N6011), .B(N8255), .C(N6006), .D(N8281));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4268 (.Y(N6023), .A(N8198), .B(N8379));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4270 (.Y(N6025), .A(N8288), .B(N8460));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4277 (.Y(N6032), .A(N4326), .B(N4822));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6178 (.Y(N6034), .A(N4262), .B(N5224), .C(N4477));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6179 (.Y(N6036), .AN(N8238), .BN(N8455), .C(N8602), .D(N6023));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6181 (.Y(N6038), .AN(N6025), .B(N8182), .C(N6032), .D(N8178));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6182 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[54]), .AN(N6038), .B(N6036), .C(N6034));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4293 (.Y(N6049), .A(N8206), .B(N8238));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4299 (.Y(N6055), .A(N6743), .B(N8521));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4306 (.Y(N6062), .A(N6809), .B(N4677));
NAND2XL hyperpropagate_3_1_A_I7515 (.Y(N8973), .A(N8539), .B(N8198));
NOR2XL hyperpropagate_3_1_A_I7516 (.Y(N6067), .A(N6833), .B(N8973));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6187 (.Y(N6068), .AN(N6055), .B(N8223), .C(N6062), .D(N8304));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6188 (.Y(N6072), .AN(N6049), .B(N8413), .C(N6067), .D(N8325));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6189 (.Y(N6070), .A(N8567), .B(N6065), .C(N5738), .D(N6068));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4315 (.Y(N6074), .A(N5156), .B(N4576));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4317 (.Y(N6073), .A(N6072), .B(N6070));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4319 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[55]), .A(N6074), .B(N6073));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4329 (.Y(N6086), .A(N8299), .B(N8439));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4339 (.Y(N6096), .A(N8260), .B(N8325));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4342 (.Y(N6102), .A(N8562), .B(N5429));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6557 (.Y(N6101), .A(N8528), .B(N8336), .C(N6753), .D(N8308));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4347 (.Y(N6104), .A(N6086), .B(N6793));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6194 (.Y(N6110), .AN(N6096), .B(N8508), .C(N6101), .D(N6727));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6196 (.Y(N6109), .A(N8467), .B(N8474), .C(N8129), .D(N6104));
NAND3XL hyperpropagate_4_1_A_I7517 (.Y(N8982), .A(N8551), .B(N8394), .C(N6102));
NOR2XL hyperpropagate_4_1_A_I7518 (.Y(N6114), .A(N6110), .B(N8982));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6198 (.Y(N6113), .A(N111), .B(N4500), .C(N4755), .D(N6109));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4358 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[56]), .A(N6114), .B(N6113));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4364 (.Y(N6121), .A(N8308), .B(N8299));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4372 (.Y(N6129), .A(N159), .B(N4500));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4378 (.Y(N6135), .A(N6142), .B(N4290));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6200 (.Y(N6138), .A(N8575), .B(N8609), .C(N6121));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6201 (.Y(N6145), .AN(N8439), .BN(N8233), .C(N6837), .D(N6139));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6204 (.Y(N6144), .AN(N8595), .B(N8496), .C(N6138), .D(N8426));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6205 (.Y(N6147), .AN(N6727), .BN(N6769), .C(N6135), .D(N6144));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6206 (.Y(N6149), .A(N8255), .B(N8521), .C(N6147));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6207 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[57]), .AN(N6149), .B(N6129), .C(N6145));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4403 (.Y(N6160), .A(N8227), .B(N8362));
NAND2XL hyperpropagate_3_1_A_I7519 (.Y(N8988), .A(N8354), .B(N8242));
NOR2XL hyperpropagate_3_1_A_I7520 (.Y(N6174), .A(N4647), .B(N8988));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4418 (.Y(N6175), .A(N6789), .B(N6809));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4419 (.Y(N6181), .A(N5128), .B(N5885));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6212 (.Y(N6178), .AN(N8188), .BN(N6769), .C(N8609), .D(N6160));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6214 (.Y(N6187), .A(N8539), .B(N8467), .C(N8299), .D(N6181));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6215 (.Y(N6183), .A(N8567), .B(N4614), .C(N6172), .D(N8595));
NAND3XL hyperpropagate_4_1_A_I7521 (.Y(N8997), .A(N8310), .B(N8521), .C(N6174));
NOR2XL hyperpropagate_4_1_A_I7522 (.Y(N6189), .A(N6183), .B(N8997));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6218 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[58]), .AN(N6187), .B(N6175), .C(N6189), .D(N6178));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4438 (.Y(N6195), .A(N8386), .B(N8202));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4446 (.Y(N6485), .A(N8535), .B(N8264));
NAND2XL hyperpropagate_3_1_A_I7523 (.Y(N9003), .A(N8486), .B(N8411));
NOR2XL hyperpropagate_3_1_A_I7524 (.Y(N6207), .A(N6485), .B(N9003));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6222 (.Y(N6213), .A(N8130), .B(N6195), .C(N6212));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6223 (.Y(N6214), .AN(N6823), .B(N8178), .C(N6207), .D(N8185));
NAND2XL hyperpropagate_3_1_A_I7525 (.Y(N9010), .A(N8242), .B(N8299));
NOR2XL hyperpropagate_3_1_A_I7526 (.Y(N6216), .A(N6142), .B(N9010));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6226 (.Y(N6218), .AN(N6213), .B(N8281), .C(N6216), .D(N8218));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6227 (.Y(N6220), .A(N6787), .B(N6214), .C(N6218));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6228 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[59]), .A(N8332), .B(N8350), .C(N8455), .D(N6220));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4473 (.Y(N6230), .A(N8426), .B(N8288));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4474 (.Y(N6231), .A(N8264), .B(N8543));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6231 (.Y(N6245), .AN(N8539), .BN(N8174), .C(N4389), .D(N5967));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6232 (.Y(N6247), .AN(N8212), .BN(N6753), .C(N6230), .D(N6231));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6558 (.Y(N6251), .A(N6212), .B(N4477), .C(N4826), .D(N6809));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6234 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[60]), .A(N6247), .B(N6245), .C(N6251));
NAND2XL hyperpropagate_3_1_A_I7527 (.Y(N9017), .A(N8435), .B(N8478));
NOR2XL hyperpropagate_3_1_A_I7528 (.Y(N6263), .A(N5148), .B(N9017));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4507 (.Y(N6264), .A(N8255), .B(N8346));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4508 (.Y(N6280), .A(N4410), .B(N6837));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6236 (.Y(N6267), .A(N8304), .B(N8332), .C(N8238));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4515 (.Y(N6272), .A(N8325), .B(N8464));
NAND3XL hyperpropagate_4_1_A_I7529 (.Y(N9026), .A(N8525), .B(N6739), .C(N6263));
NOR2XL hyperpropagate_4_1_A_I7530 (.Y(N6277), .A(N4656), .B(N9026));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6239 (.Y(N6279), .A(N6278), .B(N6805), .C(N6272));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I6559 (.Y(N6287), .AN(N6279), .B(N4832), .C(N6267), .D(N5562));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6242 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[61]), .AN(N6264), .B(N6280), .C(N6287), .D(N6277));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4540 (.Y(N6298), .A(N6715), .B(N6705));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4543 (.Y(N6301), .A(N8362), .B(N8417));
NAND2XL hyperpropagate_3_1_A_I7531 (.Y(N9032), .A(N8375), .B(N8455));
NOR2XL hyperpropagate_3_1_A_I7532 (.Y(N6303), .A(N6701), .B(N9032));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4554 (.Y(N6312), .A(N8562), .B(N5998));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4555 (.Y(N6313), .A(N6298), .B(N6312));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6245 (.Y(N6315), .AN(N8435), .BN(N8407), .C(N5657), .D(N6314));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6246 (.Y(N6317), .A(N6049), .B(N6301), .C(N6316));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6248 (.Y(N6320), .AN(N6313), .B(N8426), .C(N6303), .D(N8394));
NAND2XL hyperpropagate_3_1_A_I7533 (.Y(N9039), .A(N8332), .B(N8508));
NOR2XL hyperpropagate_3_1_A_I7534 (.Y(N6323), .A(N6320), .B(N9039));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6251 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[62]), .AN(N5779), .B(N6317), .C(N6323), .D(N6315));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4583 (.Y(N6346), .A(N5657), .B(N4319));
OR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6252 (.Y(N6345), .A(N144), .B(N8130), .C(N6344));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4591 (.Y(N6350), .A(N8525), .B(N8383));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6255 (.Y(N6361), .A(N6807), .B(N5078), .C(N6356));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6256 (.Y(N6358), .A(N8575), .B(N4789), .C(N6350), .D(N6354));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4603 (.Y(N6362), .A(N6361), .B(N6358));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6258 (.Y(N6364), .AN(N6346), .BN(N5264), .C(N6345), .D(N6362));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6259 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[63]), .A(N8332), .B(N8421), .C(N8407), .D(N6364));
NAND3XL hyperpropagate_4_1_A_I7535 (.Y(N9048), .A(N8366), .B(N8332), .C(N8346));
NOR2XL hyperpropagate_4_1_A_I7536 (.Y(N6397), .A(N6721), .B(N9048));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4623 (.Y(N6383), .A(N8413), .B(N8212));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6262 (.Y(N6389), .A(N4656), .B(N6813), .C(N6383));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6263 (.Y(N6391), .AN(N4737), .B(N6272), .C(N5261));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6266 (.Y(N6395), .AN(N6793), .B(N8372), .C(N6391), .D(N8455));
NAND3XL hyperpropagate_4_1_A_I7537 (.Y(N9056), .A(N8304), .B(N8299), .C(N6389));
NOR2XL hyperpropagate_4_1_A_I7538 (.Y(N6396), .A(N6395), .B(N9056));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4638 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[64]), .A(N6397), .B(N6396));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4657 (.Y(N6418), .A(N8547), .B(N8336));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4659 (.Y(N6420), .A(N4297), .B(N4917));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6269 (.Y(N6422), .A(N6817), .B(N4824), .C(N5423));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6560 (.Y(N6426), .AN(N8417), .BN(N8449), .C(N6695), .D(N6418));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6272 (.Y(N6429), .AN(N6801), .BN(N8605), .C(N6755), .D(N6422));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6273 (.Y(N6432), .A(N8315), .B(N8521), .C(N6426));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I5613 (.Y(N6435), .AN(N8426), .BN(N8500), .C(N6793), .D(N6432));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6275 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[65]), .AN(N6429), .B(N4365), .C(N6435), .D(N6420));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4686 (.Y(N6447), .A(N8264), .B(N8460));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4692 (.Y(N6453), .A(N5560), .B(N5791));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6279 (.Y(N6459), .AN(N5353), .B(N8397), .C(N6453), .D(N6753));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4700 (.Y(N6461), .A(N4507), .B(N5654));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6281 (.Y(N6463), .AN(N8411), .BN(N8505), .C(N4831), .D(N6447));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6282 (.Y(N6466), .A(N6350), .B(N6418), .C(N6457), .D(N6459));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6283 (.Y(N6465), .AN(N4322), .B(N8496), .C(N6461), .D(N8198));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4706 (.Y(N6467), .A(N6466), .B(N6465));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4707 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[66]), .A(N6463), .B(N6467));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6287 (.Y(N6495), .AN(N8411), .BN(N8308), .C(N4288), .D(N6485));
NAND3XL hyperpropagate_4_1_A_I7539 (.Y(N9064), .A(N8223), .B(N8354), .C(N8332));
NOR3BXL hyperpropagate_4_1_A_I10076 (.Y(N6503), .AN(N8247), .B(N9064), .C(N6195));
NAND2XL hyperpropagate_3_1_A_I7541 (.Y(N9070), .A(N8315), .B(N8474));
NOR2XL hyperpropagate_3_1_A_I7542 (.Y(N6497), .A(N6793), .B(N9070));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6292 (.Y(N6501), .A(N4762), .B(N6833), .C(N6837), .D(N5998));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6293 (.Y(N6500), .AN(N5885), .BN(N4574), .C(N6497), .D(N6495));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4741 (.Y(N6502), .A(N6501), .B(N6500));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4743 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[67]), .A(N6503), .B(N6502));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4747 (.Y(N6508), .A(N8202), .B(N8294));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4748 (.Y(N6509), .A(N8247), .B(N8174));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4750 (.Y(N6511), .A(N8407), .B(N8277));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4756 (.Y(N6517), .A(N6777), .B(N6769));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4762 (.Y(N6523), .A(N8603), .B(N5566));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6295 (.Y(N6525), .AN(N6517), .B(N8535), .C(N6509), .D(N8508));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6298 (.Y(N6539), .A(N4443), .B(N8607), .C(N6508), .D(N6301));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6299 (.Y(N6536), .AN(N4365), .BN(N6523), .C(N4537), .D(N6511));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I6301 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[68]), .AN(N6531), .BN(N6525), .C(N6539), .D(N6536));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4788 (.Y(N6549), .A(N8379), .B(N8401));
NAND2XL hyperpropagate_3_1_A_I7543 (.Y(N9077), .A(N8470), .B(N8336));
NOR2XL hyperpropagate_3_1_A_I7544 (.Y(N6558), .A(N6835), .B(N9077));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6304 (.Y(N6564), .AN(N6563), .B(N8242), .C(N8426));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6306 (.Y(N6569), .AN(N6549), .B(N8366), .C(N6558), .D(N8508));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6307 (.Y(N6568), .A(N5302), .B(N6508), .C(N6564));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6308 (.Y(N6570), .A(N6795), .B(N8579), .C(N6354), .D(N6569));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4810 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[69]), .A(N6568), .B(N6570));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4827 (.Y(N6593), .A(N6835), .B(N6813));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4828 (.Y(N6595), .A(N5768), .B(N5427));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4829 (.Y(N6591), .A(N8598), .B(N6695));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4830 (.Y(N6592), .A(N6795), .B(N8609));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I6309 (.Y(N6594), .A(N8421), .B(N8198), .C(N6593));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6312 (.Y(N6601), .AN(N6591), .BN(N6592), .C(N8579), .D(N6595));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I6313 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[70]), .AN(N6594), .B(N8379), .C(N6601), .D(N8535));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I6314 (.Y(N6624), .AN(N5595), .B(N8375), .C(N8249));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4862 (.Y(N6625), .A(N6624), .B(N6805));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4863 (.Y(N6626), .A(N6795), .B(N6811));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6316 (.Y(N6633), .A(N4897), .B(N6695), .C(N4297));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4868 (.Y(N6631), .A(N6626), .B(N6625));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I6317 (.Y(N6632), .A(N5594), .B(N6813), .C(N8609), .D(N6631));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4871 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[71]), .A(N6633), .B(N6632));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I4877 (.Y(N6640), .A(N8299), .B(N8535));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I4891 (.Y(N6654), .A(N8607), .B(N4296));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I6319 (.Y(N6656), .AN(N8508), .BN(N8383), .C(N6835), .D(N8609));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6320 (.Y(N6658), .A(N4984), .B(N6823), .C(N6640));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I6321 (.Y(N6660), .A(N4480), .B(N6809), .C(N8598));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I6561 (.Y(inst_cellmath__195__80__2WWMM_2WWMM_out0[72]), .A(N6654), .B(N6656), .C(N6660), .D(N6658));
assign inst_cellmath__195__80__2WWMM_2WWMM_out0[22] = 1'B0;
endmodule

module cynw_cm_float_sin_inst_cellmath__198_0_bdw1946085813_bdw (
	inst_cellmath__198_0_out0,
	inst_cellmath__198_0_in0,
	inst_cellmath__198_0_in1
	); /* architecture "gate_level" */ 
output [32:0] inst_cellmath__198_0_out0;
input [15:0] inst_cellmath__198_0_in0;
input [0:0] inst_cellmath__198_0_in1;
wire N102,N106,N108,N110,N112,N114,N116 
	,N118,N120,N122,N124,N126,N128,N130,N148 
	,N150,N152,N154,N156,N158,N160,N162,N164 
	,N166,N168,N170,N172,N174,N188,N192,N194 
	,N196,N198,N200,N202,N204,N206,N208,N210 
	,N212,N214,N216,N230,N234,N236,N238,N240 
	,N242,N244,N246,N248,N250,N252,N254,N256 
	,N270,N274,N276,N278,N280,N282,N284,N286 
	,N288,N290,N292,N294,N308,N312,N314,N316 
	,N318,N320,N322,N324,N326,N328,N330,N344 
	,N348,N350,N352,N354,N356,N358,N360,N362 
	,N364,N378,N382,N384,N386,N388,N390,N392 
	,N394,N396,N410,N414,N416,N418,N420,N422 
	,N424,N426,N440,N444,N446,N448,N450,N452 
	,N454,N468,N472,N474,N476,N478,N480,N494 
	,N498,N500,N502,N504,N518,N522,N524,N526 
	,N540,N544,N546,N560,N564,N578,N598,N599 
	,N600,N601,N602,N603,N604,N605,N606,N607 
	,N608,N609,N610,N611,N612,N613,N614,N615 
	,N616,N617,N618,N619,N620,N621,N622,N623 
	,N624,N625,N626,N627,N628,N629,N630,N631 
	,N632,N633,N634,N635,N636,N637,N638,N639 
	,N640,N641,N642,N643,N644,N645,N646,N647 
	,N648,N649,N650,N651,N652,N653,N654,N655 
	,N656,N657,N658,N659,N660,N661,N662,N663 
	,N664,N665,N666,N667,N668,N669,N670,N671 
	,N672,N673,N674,N675,N676,N677,N678,N679 
	,N680,N681,N682,N683,N684,N685,N686,N687 
	,N688,N689,N690,N691,N692,N693,N694,N695 
	,N696,N697,N698,N699,N700,N701,N702,N703 
	,N704,N705,N706,N707,N708,N709,N710,N711 
	,N712,N715,N716,N717,N718,N719,N720,N721 
	,N722,N723,N724,N725,N726,N727,N728,N729 
	,N730,N731,N732,N733,N734,N735,N736,N737 
	,N738,N739,N740,N741,N742,N743,N744,N745 
	,N746,N747,N748,N749,N750,N751,N752,N753 
	,N754,N755,N756,N757,N758,N759,N760,N761 
	,N762,N763,N764,N765,N766,N767,N768,N769 
	,N770,N771,N772,N773,N774,N775,N776,N777 
	,N778,N779,N780,N781,N782,N783,N784,N785 
	,N786,N787,N788,N789,N790,N791,N792,N793 
	,N794,N795,N796,N797,N798,N799,N800,N801 
	,N802,N803,N804,N805,N806,N807,N808,N809 
	,N810,N811,N812,N813,N814,N815,N816,N817 
	,N818,N819,N820,N821,N822,N823,N824,N825 
	,N826,N827,N828,N829,N830,N831,N832,N833 
	,N834,N835,N836,N837,N838,N839,N840,N841 
	,N842,N843,N844,N847,N857,N865,N877,N889 
	,N905,N921,N941,N945,N969,N971,N993,N996 
	,N999,N1002,N1005,N1008,N1011,N1014,N1017,N1029 
	,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038 
	,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046 
	,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054 
	,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062 
	,N1063,N1064,N1065,N1066,N1067,N1068,N1073,N1077 
	,N1078,N1081,N1082,N1085,N1086,N1089,N1090,N1093 
	,N1094,N1097,N1098,N1101,N1102,N1107,N1108,N1113 
	,N1114,N1117,N1118,N1123,N1124,N1147,N1149,N1150 
	,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158 
	,N1159,N1160,N1165,N1167,N1169,N1170,N1171,N1172 
	,N1173,N1174,N1175,N1176,N1185,N1187,N1189,N1191 
	,N1224,N1227,N1230,N1233,N1236,N1239,N1242,N1245 
	,N1248,N1251,N1254,N1257,N1260,N1263,N1266,N1269 
	,N1272,N1275,N1278,N1281,N1292,N1293,N1295,N1296 
	,N1298,N1299,N1301,N1302,N1304,N1305,N1307,N1308 
	,N1310,N1311,N1313,N1314,N1316,N1317,N1319,N1320 
	,N1322,N1323,N1529,N1538,N1554,N1563,N1577,N1578 
	,N1579,N1580,N1582,N1583,N1589,N1596,N1602,N1603 
	,N1609,N1616,N1618,N1626,N1627,N1632,N1633,N1638 
	,N1640,N1641,N1647,N1649,N1650,N1652,N1654,N1655 
	,N1656,N1658,N1662,N1664,N1669,N1671,N1672,N1673 
	,N1679,N1680,N1690,N1691,N1705,N1706,N1721,N1722 
	,N1746,N1747,N1754,N1755,N1766,N1767,N1774,N1775 
	,N1776,N1777,N1778,N1795,N1801;
INVX1 inst_cellmath__198_0_I931 (.Y(N1577), .A(inst_cellmath__198_0_in0[1]));
INVX2 inst_cellmath__198_0_I932 (.Y(N1578), .A(N1577));
INVXL inst_cellmath__198_0_I937 (.Y(N1583), .A(N1578));
INVX1 inst_cellmath__198_0_I936 (.Y(N1582), .A(N1578));
INVX1 inst_cellmath__198_0_I934 (.Y(N1580), .A(N1578));
INVXL inst_cellmath__198_0_I933 (.Y(N1579), .A(N1578));
INVX1 inst_cellmath__198_0_I943 (.Y(N1589), .A(inst_cellmath__198_0_in0[2]));
INVX1 inst_cellmath__198_0_I950 (.Y(N1596), .A(inst_cellmath__198_0_in0[3]));
INVXL inst_cellmath__198_0_I957 (.Y(N1603), .A(inst_cellmath__198_0_in0[4]));
INVXL inst_cellmath__198_0_I956 (.Y(N1602), .A(inst_cellmath__198_0_in0[4]));
INVX1 inst_cellmath__198_0_I963 (.Y(N1609), .A(inst_cellmath__198_0_in0[5]));
INVX1 inst_cellmath__198_0_I970 (.Y(N1616), .A(inst_cellmath__198_0_in0[6]));
INVX1 inst_cellmath__198_0_I972 (.Y(N1618), .A(inst_cellmath__198_0_in0[7]));
INVX1 inst_cellmath__198_0_I980 (.Y(N1626), .A(inst_cellmath__198_0_in0[8]));
INVX1 inst_cellmath__198_0_I981 (.Y(N1627), .A(inst_cellmath__198_0_in0[9]));
INVX1 inst_cellmath__198_0_I987 (.Y(N1633), .A(inst_cellmath__198_0_in0[10]));
INVXL inst_cellmath__198_0_I986 (.Y(N1632), .A(inst_cellmath__198_0_in0[10]));
INVXL inst_cellmath__198_0_I995 (.Y(N1641), .A(inst_cellmath__198_0_in0[11]));
INVXL inst_cellmath__198_0_I994 (.Y(N1640), .A(inst_cellmath__198_0_in0[11]));
INVXL inst_cellmath__198_0_I992 (.Y(N1638), .A(inst_cellmath__198_0_in0[11]));
INVX1 inst_cellmath__198_0_I1001 (.Y(N1647), .A(inst_cellmath__198_0_in0[12]));
INVXL inst_cellmath__198_0_I1003 (.Y(N1649), .A(inst_cellmath__198_0_in0[13]));
INVX1 inst_cellmath__198_0_I1004 (.Y(N1650), .A(N1649));
INVXL inst_cellmath__198_0_I1009 (.Y(N1655), .A(N1650));
INVX2 inst_cellmath__198_0_I1008 (.Y(N1654), .A(N1650));
INVXL inst_cellmath__198_0_I1006 (.Y(N1652), .A(N1650));
INVX1 inst_cellmath__198_0_I1010 (.Y(N1656), .A(inst_cellmath__198_0_in0[14]));
BUFX2 inst_cellmath__198_0_I1207 (.Y(N1658), .A(inst_cellmath__198_0_in0[15]));
INVX1 inst_cellmath__198_0_I1016 (.Y(N1662), .A(N1658));
INVXL inst_cellmath__198_0_I1018 (.Y(N1664), .A(inst_cellmath__198_0_in1[0]));
INVXL inst_cellmath__198_0_I1025 (.Y(N1671), .A(inst_cellmath__198_0_in0[0]));
INVXL inst_cellmath__198_0_I1023 (.Y(N1669), .A(inst_cellmath__198_0_in0[0]));
INVXL inst_cellmath__198_0_I21 (.Y(inst_cellmath__198_0_out0[0]), .A(N1671));
OR2XL inst_cellmath__198_0_I23 (.Y(N102), .A(N1669), .B(N1583));
NOR2BX1 inst_cellmath__198_0_I1173 (.Y(N826), .AN(inst_cellmath__198_0_in0[2]), .B(N1671));
NOR2XL inst_cellmath__198_0_I25 (.Y(N106), .A(N1671), .B(N1596));
NOR2XL inst_cellmath__198_0_I26 (.Y(N108), .A(N1671), .B(N1603));
NOR2BX1 inst_cellmath__198_0_I1174 (.Y(N110), .AN(inst_cellmath__198_0_in0[5]), .B(N1671));
NOR2BX1 inst_cellmath__198_0_I1175 (.Y(N112), .AN(inst_cellmath__198_0_in0[6]), .B(N1669));
NOR2XL inst_cellmath__198_0_I29 (.Y(N114), .A(N1669), .B(N1618));
NOR2XL inst_cellmath__198_0_I30 (.Y(N116), .A(N1669), .B(N1626));
NOR2XL inst_cellmath__198_0_I31 (.Y(N118), .A(N1669), .B(N1627));
NOR2BX1 inst_cellmath__198_0_I1209 (.Y(N120), .AN(inst_cellmath__198_0_in0[10]), .B(N1671));
NOR2XL inst_cellmath__198_0_I33 (.Y(N122), .A(N1671), .B(N1641));
NOR2BX1 inst_cellmath__198_0_I1248 (.Y(N124), .AN(inst_cellmath__198_0_in0[12]), .B(N1671));
NOR2XL inst_cellmath__198_0_I35 (.Y(N126), .A(N1671), .B(N1655));
NOR2XL inst_cellmath__198_0_I36 (.Y(N128), .A(N1669), .B(N1656));
NOR2BX1 inst_cellmath__198_0_I1178 (.Y(N130), .AN(N1658), .B(N1669));
OR2XL inst_cellmath__198_0_I38 (.Y(N598), .A(N1669), .B(N1664));
NOR2XL inst_cellmath__198_0_I45 (.Y(N148), .A(N1582), .B(N1589));
NOR2XL inst_cellmath__198_0_I46 (.Y(N150), .A(N1582), .B(N1596));
NOR2XL inst_cellmath__198_0_I47 (.Y(N152), .A(N1582), .B(N1602));
NOR2XL inst_cellmath__198_0_I48 (.Y(N154), .A(N1582), .B(N1609));
NOR2XL inst_cellmath__198_0_I49 (.Y(N156), .A(N1582), .B(N1616));
NOR2XL inst_cellmath__198_0_I50 (.Y(N158), .A(N1582), .B(N1618));
NOR2XL inst_cellmath__198_0_I51 (.Y(N160), .A(N1582), .B(N1626));
NOR2XL inst_cellmath__198_0_I52 (.Y(N162), .A(N1582), .B(N1627));
NOR2XL inst_cellmath__198_0_I53 (.Y(N164), .A(N1580), .B(N1633));
NOR2XL inst_cellmath__198_0_I54 (.Y(N166), .A(N1580), .B(N1640));
NOR2XL inst_cellmath__198_0_I55 (.Y(N168), .A(N1580), .B(N1647));
NOR2XL inst_cellmath__198_0_I56 (.Y(N170), .A(N1580), .B(N1654));
NOR2XL inst_cellmath__198_0_I57 (.Y(N172), .A(N1579), .B(N1656));
NOR2XL inst_cellmath__198_0_I58 (.Y(N174), .A(N1579), .B(N1662));
OR2XL inst_cellmath__198_0_I2358 (.Y(N599), .A(N1579), .B(N1664));
INVXL inst_cellmath__198_0_I64 (.Y(N188), .A(N1589));
NOR2XL inst_cellmath__198_0_I66 (.Y(N192), .A(N1589), .B(N1596));
NOR2XL inst_cellmath__198_0_I67 (.Y(N194), .A(N1589), .B(N1602));
NOR2XL inst_cellmath__198_0_I68 (.Y(N196), .A(N1589), .B(N1609));
NOR2XL inst_cellmath__198_0_I69 (.Y(N198), .A(N1589), .B(N1616));
NOR2XL inst_cellmath__198_0_I70 (.Y(N200), .A(N1589), .B(N1618));
NOR2XL inst_cellmath__198_0_I71 (.Y(N202), .A(N1589), .B(N1626));
NOR2XL inst_cellmath__198_0_I72 (.Y(N204), .A(N1589), .B(N1627));
NOR2XL inst_cellmath__198_0_I73 (.Y(N206), .A(N1589), .B(N1633));
NOR2XL inst_cellmath__198_0_I74 (.Y(N208), .A(N1589), .B(N1640));
NOR2XL inst_cellmath__198_0_I75 (.Y(N210), .A(N1589), .B(N1647));
NOR2XL inst_cellmath__198_0_I76 (.Y(N212), .A(N1589), .B(N1654));
NOR2XL inst_cellmath__198_0_I77 (.Y(N214), .A(N1589), .B(N1656));
NOR2XL inst_cellmath__198_0_I78 (.Y(N216), .A(N1589), .B(N1662));
OR2XL inst_cellmath__198_0_I79 (.Y(N600), .A(N1589), .B(N1664));
INVXL inst_cellmath__198_0_I84 (.Y(N230), .A(N1596));
NOR2XL inst_cellmath__198_0_I86 (.Y(N234), .A(N1596), .B(N1602));
NOR2XL inst_cellmath__198_0_I87 (.Y(N236), .A(N1596), .B(N1609));
NOR2XL inst_cellmath__198_0_I88 (.Y(N238), .A(N1596), .B(N1616));
NOR2XL inst_cellmath__198_0_I89 (.Y(N240), .A(N1596), .B(N1618));
NOR2XL inst_cellmath__198_0_I90 (.Y(N242), .A(N1596), .B(N1626));
NOR2XL inst_cellmath__198_0_I91 (.Y(N244), .A(N1596), .B(N1627));
NOR2XL inst_cellmath__198_0_I92 (.Y(N246), .A(N1596), .B(N1633));
NOR2XL inst_cellmath__198_0_I93 (.Y(N248), .A(N1596), .B(N1640));
NOR2XL inst_cellmath__198_0_I94 (.Y(N250), .A(N1596), .B(N1647));
NOR2XL inst_cellmath__198_0_I95 (.Y(N252), .A(N1596), .B(N1654));
NOR2XL inst_cellmath__198_0_I96 (.Y(N254), .A(N1596), .B(N1656));
NOR2XL inst_cellmath__198_0_I97 (.Y(N256), .A(N1596), .B(N1662));
OR2XL inst_cellmath__198_0_I98 (.Y(N601), .A(N1596), .B(N1664));
INVXL inst_cellmath__198_0_I103 (.Y(N270), .A(N1603));
NOR2XL inst_cellmath__198_0_I105 (.Y(N274), .A(N1603), .B(N1609));
NOR2XL inst_cellmath__198_0_I106 (.Y(N276), .A(N1603), .B(N1616));
NOR2XL inst_cellmath__198_0_I107 (.Y(N278), .A(N1602), .B(N1618));
NOR2XL inst_cellmath__198_0_I108 (.Y(N280), .A(N1602), .B(N1626));
NOR2XL inst_cellmath__198_0_I109 (.Y(N282), .A(N1602), .B(N1627));
NOR2XL inst_cellmath__198_0_I110 (.Y(N284), .A(N1602), .B(N1633));
NOR2XL inst_cellmath__198_0_I111 (.Y(N286), .A(N1603), .B(N1640));
NOR2XL inst_cellmath__198_0_I112 (.Y(N288), .A(N1603), .B(N1647));
NOR2XL inst_cellmath__198_0_I113 (.Y(N290), .A(N1603), .B(N1654));
NOR2XL inst_cellmath__198_0_I114 (.Y(N292), .A(N1603), .B(N1656));
NOR2XL inst_cellmath__198_0_I115 (.Y(N294), .A(N1602), .B(N1662));
OR2XL inst_cellmath__198_0_I116 (.Y(N602), .A(N1603), .B(N1664));
INVXL inst_cellmath__198_0_I121 (.Y(N308), .A(N1609));
NOR2XL inst_cellmath__198_0_I123 (.Y(N312), .A(N1609), .B(N1616));
NOR2XL inst_cellmath__198_0_I124 (.Y(N314), .A(N1609), .B(N1618));
NOR2XL inst_cellmath__198_0_I125 (.Y(N316), .A(N1609), .B(N1626));
NOR2XL inst_cellmath__198_0_I126 (.Y(N318), .A(N1609), .B(N1627));
NOR2XL inst_cellmath__198_0_I127 (.Y(N320), .A(N1609), .B(N1632));
NOR2XL inst_cellmath__198_0_I128 (.Y(N322), .A(N1609), .B(N1641));
NOR2XL inst_cellmath__198_0_I129 (.Y(N324), .A(N1609), .B(N1647));
NOR2XL inst_cellmath__198_0_I130 (.Y(N326), .A(N1609), .B(N1654));
NOR2XL inst_cellmath__198_0_I131 (.Y(N328), .A(N1609), .B(N1656));
NOR2XL inst_cellmath__198_0_I132 (.Y(N330), .A(N1609), .B(N1662));
OR2XL inst_cellmath__198_0_I133 (.Y(N603), .A(N1609), .B(N1664));
INVXL inst_cellmath__198_0_I138 (.Y(N344), .A(N1616));
NOR2XL inst_cellmath__198_0_I140 (.Y(N348), .A(N1616), .B(N1618));
NOR2XL inst_cellmath__198_0_I141 (.Y(N350), .A(N1616), .B(N1626));
NOR2XL inst_cellmath__198_0_I142 (.Y(N352), .A(N1616), .B(N1627));
NOR2XL inst_cellmath__198_0_I143 (.Y(N354), .A(N1616), .B(N1632));
NOR2XL inst_cellmath__198_0_I144 (.Y(N356), .A(N1616), .B(N1641));
NOR2XL inst_cellmath__198_0_I145 (.Y(N358), .A(N1616), .B(N1647));
NOR2XL inst_cellmath__198_0_I146 (.Y(N360), .A(N1616), .B(N1654));
NOR2XL inst_cellmath__198_0_I147 (.Y(N362), .A(N1616), .B(N1656));
NOR2XL inst_cellmath__198_0_I148 (.Y(N364), .A(N1616), .B(N1662));
OR2XL inst_cellmath__198_0_I149 (.Y(N604), .A(N1616), .B(N1664));
INVXL inst_cellmath__198_0_I154 (.Y(N378), .A(N1618));
NOR2XL inst_cellmath__198_0_I156 (.Y(N382), .A(N1618), .B(N1626));
NOR2XL inst_cellmath__198_0_I157 (.Y(N384), .A(N1618), .B(N1627));
NOR2XL inst_cellmath__198_0_I158 (.Y(N386), .A(N1618), .B(N1632));
NOR2XL inst_cellmath__198_0_I159 (.Y(N388), .A(N1618), .B(N1641));
NOR2XL inst_cellmath__198_0_I160 (.Y(N390), .A(N1618), .B(N1647));
NOR2XL inst_cellmath__198_0_I161 (.Y(N392), .A(N1618), .B(N1654));
NOR2XL inst_cellmath__198_0_I162 (.Y(N394), .A(N1618), .B(N1656));
NOR2XL inst_cellmath__198_0_I163 (.Y(N396), .A(N1618), .B(N1662));
OR2XL inst_cellmath__198_0_I164 (.Y(N605), .A(N1618), .B(N1664));
INVXL inst_cellmath__198_0_I169 (.Y(N410), .A(N1626));
NOR2XL inst_cellmath__198_0_I171 (.Y(N414), .A(N1626), .B(N1627));
NOR2XL inst_cellmath__198_0_I172 (.Y(N416), .A(N1626), .B(N1632));
NOR2XL inst_cellmath__198_0_I173 (.Y(N418), .A(N1626), .B(N1641));
NOR2XL inst_cellmath__198_0_I174 (.Y(N420), .A(N1626), .B(N1647));
NOR2XL inst_cellmath__198_0_I175 (.Y(N422), .A(N1626), .B(N1654));
NOR2XL inst_cellmath__198_0_I176 (.Y(N424), .A(N1626), .B(N1656));
NOR2XL inst_cellmath__198_0_I177 (.Y(N426), .A(N1626), .B(N1662));
OR2XL inst_cellmath__198_0_I178 (.Y(N606), .A(N1626), .B(N1664));
INVXL inst_cellmath__198_0_I183 (.Y(N440), .A(N1627));
NOR2XL inst_cellmath__198_0_I185 (.Y(N444), .A(N1627), .B(N1632));
NOR2XL inst_cellmath__198_0_I186 (.Y(N446), .A(N1627), .B(N1638));
NOR2XL inst_cellmath__198_0_I187 (.Y(N448), .A(N1627), .B(N1647));
NOR2XL inst_cellmath__198_0_I188 (.Y(N450), .A(N1627), .B(N1652));
NOR2XL inst_cellmath__198_0_I189 (.Y(N452), .A(N1627), .B(N1656));
NOR2XL inst_cellmath__198_0_I190 (.Y(N454), .A(N1627), .B(N1662));
OR2XL inst_cellmath__198_0_I191 (.Y(N607), .A(N1627), .B(N1664));
INVXL inst_cellmath__198_0_I196 (.Y(N468), .A(N1633));
NOR2XL inst_cellmath__198_0_I198 (.Y(N472), .A(N1633), .B(N1638));
NOR2XL inst_cellmath__198_0_I199 (.Y(N474), .A(N1633), .B(N1647));
NOR2XL inst_cellmath__198_0_I200 (.Y(N476), .A(N1632), .B(N1652));
NOR2XL inst_cellmath__198_0_I201 (.Y(N478), .A(N1632), .B(N1656));
NOR2XL inst_cellmath__198_0_I202 (.Y(N480), .A(N1632), .B(N1662));
OR2XL inst_cellmath__198_0_I203 (.Y(N608), .A(N1633), .B(N1664));
INVXL inst_cellmath__198_0_I208 (.Y(N494), .A(N1638));
NOR2XL inst_cellmath__198_0_I210 (.Y(N498), .A(N1638), .B(N1647));
NOR2XL inst_cellmath__198_0_I211 (.Y(N500), .A(N1638), .B(N1652));
NOR2XL inst_cellmath__198_0_I212 (.Y(N502), .A(N1638), .B(N1656));
NOR2XL inst_cellmath__198_0_I213 (.Y(N504), .A(N1638), .B(N1662));
OR2XL inst_cellmath__198_0_I214 (.Y(N609), .A(N1638), .B(N1664));
INVXL inst_cellmath__198_0_I219 (.Y(N518), .A(N1647));
NOR2XL inst_cellmath__198_0_I221 (.Y(N522), .A(N1647), .B(N1652));
NOR2XL inst_cellmath__198_0_I222 (.Y(N524), .A(N1647), .B(N1656));
NOR2XL inst_cellmath__198_0_I223 (.Y(N526), .A(N1647), .B(N1662));
OR2XL inst_cellmath__198_0_I224 (.Y(N610), .A(N1647), .B(N1664));
INVXL inst_cellmath__198_0_I229 (.Y(N540), .A(N1655));
NOR2XL inst_cellmath__198_0_I231 (.Y(N544), .A(N1655), .B(N1656));
NOR2XL inst_cellmath__198_0_I232 (.Y(N546), .A(N1655), .B(N1662));
OR2XL inst_cellmath__198_0_I233 (.Y(N611), .A(N1655), .B(N1664));
INVXL inst_cellmath__198_0_I238 (.Y(N560), .A(N1656));
NOR2XL inst_cellmath__198_0_I240 (.Y(N564), .A(N1656), .B(N1662));
OR2XL inst_cellmath__198_0_I241 (.Y(N612), .A(N1656), .B(N1664));
INVXL inst_cellmath__198_0_I246 (.Y(N578), .A(N1662));
ADDHX1 inst_cellmath__198_0_I269 (.CO(N614), .S(N613), .A(N188), .B(N148));
ADDHX1 inst_cellmath__198_0_I270 (.CO(N616), .S(N615), .A(N150), .B(N108));
ADDHX1 inst_cellmath__198_0_I271 (.CO(N618), .S(N617), .A(N110), .B(N192));
ADDFX1 inst_cellmath__198_0_I272 (.CO(N620), .S(N619), .A(N152), .B(N230), .CI(N616));
ADDHX1 inst_cellmath__198_0_I273 (.CO(N622), .S(N621), .A(N112), .B(N154));
ADDFX1 inst_cellmath__198_0_I274 (.CO(N624), .S(N623), .A(N618), .B(N194), .CI(N621));
ADDHX1 inst_cellmath__198_0_I275 (.CO(N626), .S(N625), .A(N196), .B(N114));
ADDFX1 inst_cellmath__198_0_I276 (.CO(N628), .S(N627), .A(N234), .B(N156), .CI(N270));
ADDFX1 inst_cellmath__198_0_I277 (.CO(N630), .S(N629), .A(N625), .B(N622), .CI(N624));
ADDHX1 inst_cellmath__198_0_I278 (.CO(N632), .S(N631), .A(N198), .B(N158));
ADDFX1 inst_cellmath__198_0_I279 (.CO(N634), .S(N633), .A(N116), .B(N236), .CI(N626));
ADDFX1 inst_cellmath__198_0_I280 (.CO(N636), .S(N635), .A(N628), .B(N631), .CI(N633));
ADDHX1 inst_cellmath__198_0_I281 (.CO(N638), .S(N637), .A(N308), .B(N200));
ADDFX1 inst_cellmath__198_0_I282 (.CO(N640), .S(N639), .A(N118), .B(N238), .CI(N274));
ADDFX1 inst_cellmath__198_0_I283 (.CO(N642), .S(N641), .A(N632), .B(N160), .CI(N637));
ADDFX1 inst_cellmath__198_0_I284 (.CO(N644), .S(N643), .A(N639), .B(N634), .CI(N641));
ADDHX1 inst_cellmath__198_0_I285 (.CO(N646), .S(N645), .A(N120), .B(N240));
ADDFX1 inst_cellmath__198_0_I286 (.CO(N648), .S(N647), .A(N202), .B(N162), .CI(N276));
ADDFX1 inst_cellmath__198_0_I287 (.CO(N650), .S(N649), .A(N645), .B(N638), .CI(N640));
ADDFX1 inst_cellmath__198_0_I288 (.CO(N652), .S(N651), .A(N647), .B(N642), .CI(N649));
ADDHX1 inst_cellmath__198_0_I289 (.CO(N654), .S(N653), .A(N344), .B(N312));
ADDFX1 inst_cellmath__198_0_I290 (.CO(N656), .S(N655), .A(N164), .B(N122), .CI(N204));
ADDFX1 inst_cellmath__198_0_I291 (.CO(N658), .S(N657), .A(N278), .B(N242), .CI(N653));
ADDFX1 inst_cellmath__198_0_I292 (.CO(N660), .S(N659), .A(N648), .B(N646), .CI(N655));
ADDFHXL inst_cellmath__198_0_I293 (.CO(N662), .S(N661), .A(N650), .B(N657), .CI(N659));
ADDHX1 inst_cellmath__198_0_I294 (.CO(N664), .S(N663), .A(N206), .B(N314));
ADDFX1 inst_cellmath__198_0_I295 (.CO(N666), .S(N665), .A(N124), .B(N166), .CI(N244));
ADDFX1 inst_cellmath__198_0_I296 (.CO(N668), .S(N667), .A(N654), .B(N280), .CI(N663));
ADDFX1 inst_cellmath__198_0_I297 (.CO(N670), .S(N669), .A(N665), .B(N656), .CI(N658));
ADDFX1 inst_cellmath__198_0_I298 (.CO(N672), .S(N671), .A(N660), .B(N667), .CI(N669));
ADDHX1 inst_cellmath__198_0_I299 (.CO(N674), .S(N673), .A(N208), .B(N378));
ADDFX1 inst_cellmath__198_0_I300 (.CO(N676), .S(N675), .A(N168), .B(N126), .CI(N348));
ADDFX1 inst_cellmath__198_0_I301 (.CO(N678), .S(N677), .A(N316), .B(N246), .CI(N282));
ADDFX1 inst_cellmath__198_0_I302 (.CO(N680), .S(N679), .A(N673), .B(N664), .CI(N666));
ADDFX1 inst_cellmath__198_0_I303 (.CO(N682), .S(N681), .A(N668), .B(N675), .CI(N677));
ADDFX1 inst_cellmath__198_0_I304 (.CO(N684), .S(N683), .A(N670), .B(N679), .CI(N681));
ADDHX1 inst_cellmath__198_0_I305 (.CO(N686), .S(N685), .A(N170), .B(N128));
ADDFX1 inst_cellmath__198_0_I306 (.CO(N688), .S(N687), .A(N248), .B(N210), .CI(N284));
ADDFX1 inst_cellmath__198_0_I307 (.CO(N690), .S(N689), .A(N350), .B(N318), .CI(N674));
ADDFX1 inst_cellmath__198_0_I308 (.CO(N692), .S(N691), .A(N676), .B(N685), .CI(N678));
ADDFX1 inst_cellmath__198_0_I309 (.CO(N694), .S(N693), .A(N687), .B(N689), .CI(N680));
ADDFX1 inst_cellmath__198_0_I310 (.CO(N696), .S(N695), .A(N682), .B(N691), .CI(N693));
ADDHX1 inst_cellmath__198_0_I311 (.CO(N698), .S(N697), .A(N212), .B(N320));
ADDFX1 inst_cellmath__198_0_I312 (.CO(N700), .S(N699), .A(N172), .B(N130), .CI(N250));
ADDFX1 inst_cellmath__198_0_I313 (.CO(N702), .S(N701), .A(N382), .B(N352), .CI(N286));
ADDFX1 inst_cellmath__198_0_I314 (.CO(N704), .S(N703), .A(N686), .B(N410), .CI(N697));
ADDFX1 inst_cellmath__198_0_I315 (.CO(N706), .S(N705), .A(N690), .B(N688), .CI(N699));
ADDFX1 inst_cellmath__198_0_I316 (.CO(N708), .S(N707), .A(N703), .B(N701), .CI(N692));
ADDFX1 inst_cellmath__198_0_I317 (.CO(N710), .S(N709), .A(N705), .B(N694), .CI(N707));
XNOR2X1 hap1_A_I898 (.Y(N711), .A(N354), .B(N174));
OR2XL hap1_A_I899 (.Y(N712), .A(N354), .B(N174));
ADDFX1 inst_cellmath__198_0_I319 (.CO(N716), .S(N715), .A(N252), .B(N214), .CI(N322));
ADDFX1 inst_cellmath__198_0_I320 (.CO(N718), .S(N717), .A(N598), .B(N288), .CI(N384));
ADDFX1 inst_cellmath__198_0_I321 (.CO(N720), .S(N719), .A(N711), .B(N698), .CI(N700));
ADDFX1 inst_cellmath__198_0_I322 (.CO(N722), .S(N721), .A(N715), .B(N702), .CI(N704));
ADDFXL inst_cellmath__198_0_I323 (.CO(N724), .S(N723), .A(N719), .B(N717), .CI(N706));
ADDFHXL inst_cellmath__198_0_I324 (.CO(N726), .S(N725), .A(N708), .B(N721), .CI(N723));
ADDFX1 inst_cellmath__198_0_I325 (.CO(N728), .S(N727), .A(N324), .B(N356), .CI(N216));
ADDFX1 inst_cellmath__198_0_I326 (.CO(N730), .S(N729), .A(N414), .B(N386), .CI(N254));
ADDFX1 inst_cellmath__198_0_I327 (.CO(N732), .S(N731), .A(N599), .B(N440), .CI(N290));
ADDFX1 inst_cellmath__198_0_I328 (.CO(N734), .S(N733), .A(N716), .B(N712), .CI(N718));
ADDFX1 inst_cellmath__198_0_I329 (.CO(N736), .S(N735), .A(N731), .B(N727), .CI(N729));
ADDFXL inst_cellmath__198_0_I330 (.CO(N738), .S(N737), .A(N722), .B(N720), .CI(N733));
ADDFXL inst_cellmath__198_0_I331 (.CO(N740), .S(N739), .A(N724), .B(N735), .CI(N737));
ADDFX1 inst_cellmath__198_0_I332 (.CO(N742), .S(N741), .A(N326), .B(N358), .CI(N388));
ADDFX1 inst_cellmath__198_0_I333 (.CO(N744), .S(N743), .A(N600), .B(N256), .CI(N292));
ADDFXL inst_cellmath__198_0_I334 (.CO(N746), .S(N745), .A(N728), .B(N416), .CI(N732));
ADDFX1 inst_cellmath__198_0_I335 (.CO(N748), .S(N747), .A(N741), .B(N730), .CI(N743));
ADDFXL inst_cellmath__198_0_I336 (.CO(N750), .S(N749), .A(N745), .B(N734), .CI(N736));
ADDFXL inst_cellmath__198_0_I337 (.CO(N752), .S(N751), .A(N738), .B(N747), .CI(N749));
ADDFX1 inst_cellmath__198_0_I338 (.CO(N754), .S(N753), .A(N360), .B(N468), .CI(N328));
ADDFX1 inst_cellmath__198_0_I339 (.CO(N756), .S(N755), .A(N444), .B(N390), .CI(N418));
ADDFX1 inst_cellmath__198_0_I340 (.CO(N758), .S(N757), .A(N601), .B(N294), .CI(N742));
ADDFX1 inst_cellmath__198_0_I341 (.CO(N760), .S(N759), .A(N753), .B(N744), .CI(N755));
ADDFX1 inst_cellmath__198_0_I342 (.CO(N762), .S(N761), .A(N757), .B(N746), .CI(N748));
ADDFX1 inst_cellmath__198_0_I343 (.CO(N764), .S(N763), .A(N750), .B(N759), .CI(N761));
ADDFX1 inst_cellmath__198_0_I344 (.CO(N766), .S(N765), .A(N330), .B(N362), .CI(N392));
ADDFX1 inst_cellmath__198_0_I345 (.CO(N768), .S(N767), .A(N420), .B(N446), .CI(N602));
ADDFX1 inst_cellmath__198_0_I346 (.CO(N770), .S(N769), .A(N756), .B(N754), .CI(N765));
ADDFX1 inst_cellmath__198_0_I347 (.CO(N772), .S(N771), .A(N758), .B(N767), .CI(N760));
ADDFX1 inst_cellmath__198_0_I348 (.CO(N774), .S(N773), .A(N762), .B(N769), .CI(N771));
ADDFX1 inst_cellmath__198_0_I349 (.CO(N776), .S(N775), .A(N472), .B(N494), .CI(N364));
ADDFX1 inst_cellmath__198_0_I350 (.CO(N778), .S(N777), .A(N603), .B(N394), .CI(N422));
ADDFX1 inst_cellmath__198_0_I351 (.CO(N780), .S(N779), .A(N766), .B(N448), .CI(N775));
ADDFX1 inst_cellmath__198_0_I352 (.CO(N782), .S(N781), .A(N777), .B(N768), .CI(N770));
ADDFX1 inst_cellmath__198_0_I353 (.CO(N784), .S(N783), .A(N772), .B(N779), .CI(N781));
ADDFX1 inst_cellmath__198_0_I354 (.CO(N786), .S(N785), .A(N396), .B(N474), .CI(N604));
ADDFX1 inst_cellmath__198_0_I355 (.CO(N788), .S(N787), .A(N424), .B(N450), .CI(N776));
ADDFX1 inst_cellmath__198_0_I356 (.CO(N790), .S(N789), .A(N785), .B(N778), .CI(N787));
ADDFX1 inst_cellmath__198_0_I357 (.CO(N792), .S(N791), .A(N782), .B(N780), .CI(N789));
ADDFX1 inst_cellmath__198_0_I358 (.CO(N794), .S(N793), .A(N518), .B(N476), .CI(N498));
ADDFX1 inst_cellmath__198_0_I359 (.CO(N796), .S(N795), .A(N605), .B(N452), .CI(N426));
ADDFX1 inst_cellmath__198_0_I360 (.CO(N798), .S(N797), .A(N793), .B(N786), .CI(N788));
ADDFX1 inst_cellmath__198_0_I361 (.CO(N800), .S(N799), .A(N797), .B(N795), .CI(N790));
ADDFX1 inst_cellmath__198_0_I362 (.CO(N802), .S(N801), .A(N478), .B(N500), .CI(N454));
ADDFX1 inst_cellmath__198_0_I363 (.CO(N804), .S(N803), .A(N794), .B(N606), .CI(N796));
ADDFX1 inst_cellmath__198_0_I364 (.CO(N806), .S(N805), .A(N798), .B(N801), .CI(N803));
ADDFX1 inst_cellmath__198_0_I365 (.CO(N808), .S(N807), .A(N480), .B(N540), .CI(N522));
ADDFX1 inst_cellmath__198_0_I366 (.CO(N810), .S(N809), .A(N607), .B(N502), .CI(N802));
ADDFX1 inst_cellmath__198_0_I367 (.CO(N812), .S(N811), .A(N804), .B(N807), .CI(N809));
ADDFX1 inst_cellmath__198_0_I368 (.CO(N814), .S(N813), .A(N524), .B(N504), .CI(N608));
ADDFX1 inst_cellmath__198_0_I369 (.CO(N816), .S(N815), .A(N813), .B(N808), .CI(N810));
ADDFX1 inst_cellmath__198_0_I370 (.CO(N818), .S(N817), .A(N526), .B(N560), .CI(N544));
ADDFX1 inst_cellmath__198_0_I371 (.CO(N820), .S(N819), .A(N814), .B(N609), .CI(N817));
ADDFX1 inst_cellmath__198_0_I372 (.CO(N822), .S(N821), .A(N610), .B(N546), .CI(N818));
ADDFX1 inst_cellmath__198_0_I373 (.CO(N824), .S(N823), .A(N564), .B(N578), .CI(N611));
NOR2XL inst_cellmath__198_0_I374 (.Y(N825), .A(N1579), .B(N102));
NOR2XL inst_cellmath__198_0_I376 (.Y(N827), .A(N106), .B(N613));
NAND2XL inst_cellmath__198_0_I377 (.Y(N828), .A(N106), .B(N613));
NOR2XL inst_cellmath__198_0_I378 (.Y(N829), .A(N614), .B(N615));
NAND2XL inst_cellmath__198_0_I379 (.Y(N830), .A(N614), .B(N615));
NOR2XL inst_cellmath__198_0_I380 (.Y(N831), .A(N617), .B(N619));
NAND2XL inst_cellmath__198_0_I381 (.Y(N832), .A(N617), .B(N619));
NOR2XL inst_cellmath__198_0_I382 (.Y(N833), .A(N620), .B(N623));
NAND2XL inst_cellmath__198_0_I383 (.Y(N834), .A(N620), .B(N623));
NOR2XL inst_cellmath__198_0_I384 (.Y(N835), .A(N627), .B(N629));
NAND2X1 inst_cellmath__198_0_I385 (.Y(N836), .A(N627), .B(N629));
NOR2XL inst_cellmath__198_0_I386 (.Y(N837), .A(N630), .B(N635));
NAND2XL inst_cellmath__198_0_I387 (.Y(N838), .A(N630), .B(N635));
NOR2XL inst_cellmath__198_0_I388 (.Y(N839), .A(N636), .B(N643));
NAND2XL inst_cellmath__198_0_I389 (.Y(N840), .A(N636), .B(N643));
NOR2XL inst_cellmath__198_0_I390 (.Y(N841), .A(N644), .B(N651));
NAND2XL inst_cellmath__198_0_I391 (.Y(N842), .A(N644), .B(N651));
NOR2XL inst_cellmath__198_0_I392 (.Y(N843), .A(N652), .B(N661));
NAND2X1 inst_cellmath__198_0_I393 (.Y(N844), .A(N652), .B(N661));
AND2XL inst_cellmath__198_0_I396 (.Y(N847), .A(N826), .B(N825));
INVXL inst_cellmath__198_0_I1026 (.Y(N1672), .A(N827));
INVXL inst_cellmath__198_0_I1027 (.Y(N1673), .A(N828));
OAI21XL inst_cellmath__198_0_I404 (.Y(N857), .A0(N1673), .A1(N847), .B0(N1672));
AOI21XL inst_cellmath__198_0_I412 (.Y(N865), .A0(N830), .A1(N857), .B0(N829));
INVXL inst_cellmath__198_0_I1033 (.Y(N1679), .A(N831));
INVXL inst_cellmath__198_0_I1034 (.Y(N1680), .A(N832));
OAI21XL inst_cellmath__198_0_I424 (.Y(N877), .A0(N1680), .A1(N865), .B0(N1679));
AOI21X1 inst_cellmath__198_0_I436 (.Y(N889), .A0(N834), .A1(N877), .B0(N833));
INVXL inst_cellmath__198_0_I1044 (.Y(N1690), .A(N835));
INVXL inst_cellmath__198_0_I1045 (.Y(N1691), .A(N836));
OAI21X2 inst_cellmath__198_0_I452 (.Y(N905), .A0(N1691), .A1(N889), .B0(N1690));
AOI21X2 inst_cellmath__198_0_I468 (.Y(N921), .A0(N838), .A1(N905), .B0(N837));
INVXL inst_cellmath__198_0_I1059 (.Y(N1705), .A(N839));
INVXL inst_cellmath__198_0_I1060 (.Y(N1706), .A(N840));
OAI21X2 inst_cellmath__198_0_I488 (.Y(N941), .A0(N1706), .A1(N921), .B0(N1705));
AOI21XL inst_cellmath__198_0_I492 (.Y(N945), .A0(N844), .A1(N841), .B0(N843));
INVXL inst_cellmath__198_0_I1075 (.Y(N1721), .A(N945));
CLKAND2X2 inst_cellmath__198_0_I1180 (.Y(N1722), .A(N844), .B(N842));
AOI21XL inst_cellmath__198_0_I516 (.Y(N969), .A0(N842), .A1(N941), .B0(N841));
AOI21X2 inst_cellmath__198_0_I518 (.Y(N971), .A0(N1722), .A1(N941), .B0(N1721));
NAND2BXL inst_cellmath__198_0_I538 (.Y(N993), .AN(N827), .B(N828));
NAND2BXL inst_cellmath__198_0_I541 (.Y(N996), .AN(N829), .B(N830));
NAND2BXL inst_cellmath__198_0_I544 (.Y(N999), .AN(N831), .B(N832));
NAND2BXL inst_cellmath__198_0_I547 (.Y(N1002), .AN(N833), .B(N834));
NAND2BXL inst_cellmath__198_0_I550 (.Y(N1005), .AN(N835), .B(N836));
NAND2BXL inst_cellmath__198_0_I553 (.Y(N1008), .AN(N837), .B(N838));
NAND2BXL inst_cellmath__198_0_I556 (.Y(N1011), .AN(N839), .B(N840));
NAND2BXL inst_cellmath__198_0_I559 (.Y(N1014), .AN(N841), .B(N842));
NAND2BXL inst_cellmath__198_0_I562 (.Y(N1017), .AN(N843), .B(N844));
XOR2XL inst_cellmath__198_0_I563 (.Y(inst_cellmath__198_0_out0[2]), .A(N1583), .B(N102));
XOR2XL inst_cellmath__198_0_I1182 (.Y(inst_cellmath__198_0_out0[3]), .A(N825), .B(N826));
XNOR2X1 inst_cellmath__198_0_I565 (.Y(inst_cellmath__198_0_out0[4]), .A(N847), .B(N993));
XOR2XL inst_cellmath__198_0_I1183 (.Y(inst_cellmath__198_0_out0[5]), .A(N857), .B(N996));
XNOR2X1 inst_cellmath__198_0_I567 (.Y(inst_cellmath__198_0_out0[6]), .A(N865), .B(N999));
XOR2XL inst_cellmath__198_0_I1184 (.Y(inst_cellmath__198_0_out0[7]), .A(N877), .B(N1002));
XNOR2X1 inst_cellmath__198_0_I569 (.Y(inst_cellmath__198_0_out0[8]), .A(N889), .B(N1005));
XOR2XL inst_cellmath__198_0_I1185 (.Y(inst_cellmath__198_0_out0[9]), .A(N905), .B(N1008));
XNOR2X1 inst_cellmath__198_0_I571 (.Y(inst_cellmath__198_0_out0[10]), .A(N921), .B(N1011));
XOR2XL inst_cellmath__198_0_I1186 (.Y(inst_cellmath__198_0_out0[11]), .A(N941), .B(N1014));
XNOR2X1 inst_cellmath__198_0_I573 (.Y(inst_cellmath__198_0_out0[12]), .A(N969), .B(N1017));
INVX2 inst_cellmath__198_0_I574 (.Y(N1029), .A(N971));
NOR2XL inst_cellmath__198_0_I575 (.Y(N1031), .A(N662), .B(N671));
NAND2XL inst_cellmath__198_0_I576 (.Y(N1032), .A(N662), .B(N671));
NOR2XL inst_cellmath__198_0_I577 (.Y(N1033), .A(N672), .B(N683));
NAND2XL inst_cellmath__198_0_I578 (.Y(N1034), .A(N672), .B(N683));
NOR2XL inst_cellmath__198_0_I579 (.Y(N1035), .A(N684), .B(N695));
NAND2XL inst_cellmath__198_0_I580 (.Y(N1036), .A(N684), .B(N695));
NOR2X1 inst_cellmath__198_0_I581 (.Y(N1037), .A(N696), .B(N709));
NAND2X1 inst_cellmath__198_0_I582 (.Y(N1038), .A(N696), .B(N709));
NOR2X1 inst_cellmath__198_0_I583 (.Y(N1039), .A(N710), .B(N725));
NAND2X4 inst_cellmath__198_0_I584 (.Y(N1040), .A(N710), .B(N725));
NOR2XL inst_cellmath__198_0_I585 (.Y(N1041), .A(N726), .B(N739));
NAND2X1 inst_cellmath__198_0_I586 (.Y(N1042), .A(N726), .B(N739));
NOR2XL inst_cellmath__198_0_I587 (.Y(N1043), .A(N740), .B(N751));
NAND2X2 inst_cellmath__198_0_I588 (.Y(N1044), .A(N740), .B(N751));
NOR2X1 inst_cellmath__198_0_I589 (.Y(N1045), .A(N752), .B(N763));
NAND2X2 inst_cellmath__198_0_I590 (.Y(N1046), .A(N752), .B(N763));
NOR2XL inst_cellmath__198_0_I591 (.Y(N1047), .A(N764), .B(N773));
NAND2X4 inst_cellmath__198_0_I592 (.Y(N1048), .A(N764), .B(N773));
NOR2XL inst_cellmath__198_0_I593 (.Y(N1049), .A(N774), .B(N783));
NAND2XL inst_cellmath__198_0_I594 (.Y(N1050), .A(N774), .B(N783));
NOR2XL inst_cellmath__198_0_I595 (.Y(N1051), .A(N784), .B(N791));
NAND2X1 inst_cellmath__198_0_I596 (.Y(N1052), .A(N784), .B(N791));
NOR2X1 inst_cellmath__198_0_I597 (.Y(N1053), .A(N792), .B(N799));
NAND2XL inst_cellmath__198_0_I598 (.Y(N1054), .A(N792), .B(N799));
NOR2XL inst_cellmath__198_0_I599 (.Y(N1055), .A(N800), .B(N805));
NAND2XL inst_cellmath__198_0_I600 (.Y(N1056), .A(N800), .B(N805));
NOR2XL inst_cellmath__198_0_I601 (.Y(N1057), .A(N806), .B(N811));
NAND2XL inst_cellmath__198_0_I602 (.Y(N1058), .A(N806), .B(N811));
NOR2XL inst_cellmath__198_0_I603 (.Y(N1059), .A(N812), .B(N815));
NAND2XL inst_cellmath__198_0_I604 (.Y(N1060), .A(N812), .B(N815));
NOR2XL inst_cellmath__198_0_I605 (.Y(N1061), .A(N816), .B(N819));
NAND2XL inst_cellmath__198_0_I606 (.Y(N1062), .A(N816), .B(N819));
NOR2XL inst_cellmath__198_0_I607 (.Y(N1063), .A(N821), .B(N820));
NAND2XL inst_cellmath__198_0_I608 (.Y(N1064), .A(N821), .B(N820));
NOR2XL inst_cellmath__198_0_I609 (.Y(N1065), .A(N823), .B(N822));
NAND2XL inst_cellmath__198_0_I610 (.Y(N1066), .A(N823), .B(N822));
NOR2XL inst_cellmath__198_0_I611 (.Y(N1067), .A(N612), .B(N824));
NAND2XL inst_cellmath__198_0_I612 (.Y(N1068), .A(N612), .B(N824));
AOI21X2 inst_cellmath__198_0_I617 (.Y(N1073), .A0(N1032), .A1(N1029), .B0(N1031));
AOI21X1 inst_cellmath__198_0_I621 (.Y(N1077), .A0(N1036), .A1(N1033), .B0(N1035));
NAND2XL inst_cellmath__198_0_I622 (.Y(N1078), .A(N1036), .B(N1034));
AOI21X4 inst_cellmath__198_0_I625 (.Y(N1081), .A0(N1040), .A1(N1037), .B0(N1039));
NAND2X4 inst_cellmath__198_0_I626 (.Y(N1082), .A(N1040), .B(N1038));
AOI21X2 inst_cellmath__198_0_I629 (.Y(N1085), .A0(N1044), .A1(N1041), .B0(N1043));
NAND2X1 inst_cellmath__198_0_I630 (.Y(N1086), .A(N1044), .B(N1042));
AOI21X2 inst_cellmath__198_0_I633 (.Y(N1089), .A0(N1048), .A1(N1045), .B0(N1047));
NAND2X2 inst_cellmath__198_0_I634 (.Y(N1090), .A(N1048), .B(N1046));
AOI21XL inst_cellmath__198_0_I637 (.Y(N1093), .A0(N1052), .A1(N1049), .B0(N1051));
NAND2XL inst_cellmath__198_0_I638 (.Y(N1094), .A(N1052), .B(N1050));
AOI21XL inst_cellmath__198_0_I641 (.Y(N1097), .A0(N1056), .A1(N1053), .B0(N1055));
NAND2XL inst_cellmath__198_0_I642 (.Y(N1098), .A(N1056), .B(N1054));
INVXL inst_cellmath__198_0_I1100 (.Y(N1746), .A(N1057));
INVXL inst_cellmath__198_0_I1101 (.Y(N1747), .A(N1058));
AOI21XL inst_cellmath__198_0_I645 (.Y(N1101), .A0(N1060), .A1(N1057), .B0(N1059));
NAND2XL inst_cellmath__198_0_I646 (.Y(N1102), .A(N1060), .B(N1058));
OAI21XL inst_cellmath__198_0_I651 (.Y(N1107), .A0(N1747), .A1(N1097), .B0(N1746));
NOR2XL inst_cellmath__198_0_I652 (.Y(N1108), .A(N1747), .B(N1098));
AOI21XL inst_cellmath__198_0_I657 (.Y(N1113), .A0(N1064), .A1(N1061), .B0(N1063));
NAND2XL inst_cellmath__198_0_I658 (.Y(N1114), .A(N1064), .B(N1062));
INVXL inst_cellmath__198_0_I1108 (.Y(N1754), .A(N1065));
INVXL inst_cellmath__198_0_I1109 (.Y(N1755), .A(N1066));
AOI21XL inst_cellmath__198_0_I661 (.Y(N1117), .A0(N1068), .A1(N1065), .B0(N1067));
NAND2XL inst_cellmath__198_0_I662 (.Y(N1118), .A(N1068), .B(N1066));
OAI21XL inst_cellmath__198_0_I667 (.Y(N1123), .A0(N1755), .A1(N1113), .B0(N1754));
NOR2XL inst_cellmath__198_0_I668 (.Y(N1124), .A(N1755), .B(N1114));
OA21X1 inst_cellmath__198_0_I1188 (.Y(N1766), .A0(N1102), .A1(N1097), .B0(N1101));
OR2XL inst_cellmath__198_0_I1189 (.Y(N1767), .A(N1102), .B(N1098));
OA21X1 inst_cellmath__198_0_I1190 (.Y(N1774), .A0(N1118), .A1(N1113), .B0(N1117));
OR2XL inst_cellmath__198_0_I1191 (.Y(N1775), .A(N1118), .B(N1114));
INVXL inst_cellmath__198_0_I1130 (.Y(N1776), .A(N1073));
OAI21X1 inst_cellmath__198_0_I691 (.Y(N1147), .A0(N1078), .A1(N1073), .B0(N1077));
OAI21X2 inst_cellmath__198_0_I693 (.Y(N1149), .A0(N1082), .A1(N1077), .B0(N1081));
NOR2X1 inst_cellmath__198_0_I694 (.Y(N1150), .A(N1082), .B(N1078));
OAI21X1 inst_cellmath__198_0_I695 (.Y(N1151), .A0(N1086), .A1(N1081), .B0(N1085));
NOR2XL inst_cellmath__198_0_I696 (.Y(N1152), .A(N1086), .B(N1082));
OAI21X1 inst_cellmath__198_0_I697 (.Y(N1153), .A0(N1090), .A1(N1085), .B0(N1089));
NOR2XL inst_cellmath__198_0_I698 (.Y(N1154), .A(N1090), .B(N1086));
OAI21XL inst_cellmath__198_0_I699 (.Y(N1155), .A0(N1094), .A1(N1089), .B0(N1093));
NOR2XL inst_cellmath__198_0_I700 (.Y(N1156), .A(N1094), .B(N1090));
OAI21XL inst_cellmath__198_0_I701 (.Y(N1157), .A0(N1767), .A1(N1093), .B0(N1766));
NOR2XL inst_cellmath__198_0_I702 (.Y(N1158), .A(N1767), .B(N1094));
OAI21XL inst_cellmath__198_0_I703 (.Y(N1159), .A0(N1775), .A1(N1766), .B0(N1774));
NOR2XL inst_cellmath__198_0_I704 (.Y(N1160), .A(N1775), .B(N1767));
INVXL inst_cellmath__198_0_I1131 (.Y(N1777), .A(N1776));
INVXL inst_cellmath__198_0_I1132 (.Y(N1778), .A(N1147));
AOI21X1 inst_cellmath__198_0_I709 (.Y(N1165), .A0(N1150), .A1(N1776), .B0(N1149));
AOI21X1 inst_cellmath__198_0_I711 (.Y(N1167), .A0(N1152), .A1(N1147), .B0(N1151));
AOI21XL inst_cellmath__198_0_I713 (.Y(N1169), .A0(N1154), .A1(N1149), .B0(N1153));
NAND2XL inst_cellmath__198_0_I714 (.Y(N1170), .A(N1154), .B(N1150));
AOI21X1 inst_cellmath__198_0_I715 (.Y(N1171), .A0(N1156), .A1(N1151), .B0(N1155));
NAND2XL inst_cellmath__198_0_I716 (.Y(N1172), .A(N1156), .B(N1152));
AOI21XL inst_cellmath__198_0_I717 (.Y(N1173), .A0(N1158), .A1(N1153), .B0(N1157));
NAND2XL inst_cellmath__198_0_I718 (.Y(N1174), .A(N1158), .B(N1154));
AOI21XL inst_cellmath__198_0_I719 (.Y(N1175), .A0(N1160), .A1(N1155), .B0(N1159));
NAND2XL inst_cellmath__198_0_I720 (.Y(N1176), .A(N1160), .B(N1156));
OAI21XL inst_cellmath__198_0_I729 (.Y(N1185), .A0(N1170), .A1(N1777), .B0(N1169));
OAI21X2 inst_cellmath__198_0_I731 (.Y(N1187), .A0(N1172), .A1(N1778), .B0(N1171));
OAI21X1 inst_cellmath__198_0_I733 (.Y(N1189), .A0(N1174), .A1(N1165), .B0(N1173));
OAI21XL inst_cellmath__198_0_I735 (.Y(N1191), .A0(N1176), .A1(N1167), .B0(N1175));
INVXL inst_cellmath__198_0_I1149 (.Y(N1795), .A(N1097));
INVXL inst_cellmath__198_0_I1155 (.Y(N1801), .A(N1113));
NAND2BXL inst_cellmath__198_0_I768 (.Y(N1224), .AN(N1031), .B(N1032));
NAND2BXL inst_cellmath__198_0_I771 (.Y(N1227), .AN(N1033), .B(N1034));
NAND2BXL inst_cellmath__198_0_I774 (.Y(N1230), .AN(N1035), .B(N1036));
NAND2BXL inst_cellmath__198_0_I777 (.Y(N1233), .AN(N1037), .B(N1038));
NAND2BXL inst_cellmath__198_0_I1194 (.Y(N1236), .AN(N1039), .B(N1040));
NAND2BXL inst_cellmath__198_0_I783 (.Y(N1239), .AN(N1041), .B(N1042));
NAND2BXL inst_cellmath__198_0_I786 (.Y(N1242), .AN(N1043), .B(N1044));
NAND2BXL inst_cellmath__198_0_I789 (.Y(N1245), .AN(N1045), .B(N1046));
NAND2BXL inst_cellmath__198_0_I792 (.Y(N1248), .AN(N1047), .B(N1048));
NAND2BXL inst_cellmath__198_0_I795 (.Y(N1251), .AN(N1049), .B(N1050));
NAND2BXL inst_cellmath__198_0_I798 (.Y(N1254), .AN(N1051), .B(N1052));
NAND2BXL inst_cellmath__198_0_I801 (.Y(N1257), .AN(N1053), .B(N1054));
NAND2BXL inst_cellmath__198_0_I804 (.Y(N1260), .AN(N1055), .B(N1056));
NAND2BXL inst_cellmath__198_0_I807 (.Y(N1263), .AN(N1057), .B(N1058));
NAND2BXL inst_cellmath__198_0_I810 (.Y(N1266), .AN(N1059), .B(N1060));
NAND2BXL inst_cellmath__198_0_I813 (.Y(N1269), .AN(N1061), .B(N1062));
NAND2BXL inst_cellmath__198_0_I816 (.Y(N1272), .AN(N1063), .B(N1064));
NAND2BXL inst_cellmath__198_0_I819 (.Y(N1275), .AN(N1065), .B(N1066));
NAND2BXL inst_cellmath__198_0_I822 (.Y(N1278), .AN(N1067), .B(N1068));
NOR2BX1 inst_cellmath__198_0_I1227 (.Y(N1281), .AN(N1662), .B(N1664));
XOR2XL inst_cellmath__198_0_I1196 (.Y(inst_cellmath__198_0_out0[13]), .A(N1029), .B(N1224));
XNOR2X1 inst_cellmath__198_0_I828 (.Y(inst_cellmath__198_0_out0[14]), .A(N1777), .B(N1227));
XNOR2X1 inst_cellmath__198_0_I829 (.Y(inst_cellmath__198_0_out0[16]), .A(N1778), .B(N1233));
XNOR2X1 inst_cellmath__198_0_I830 (.Y(inst_cellmath__198_0_out0[18]), .A(N1165), .B(N1239));
XNOR2X1 inst_cellmath__198_0_I831 (.Y(inst_cellmath__198_0_out0[20]), .A(N1167), .B(N1245));
XOR2XL inst_cellmath__198_0_I832 (.Y(inst_cellmath__198_0_out0[22]), .A(N1185), .B(N1251));
XOR2XL inst_cellmath__198_0_I833 (.Y(inst_cellmath__198_0_out0[24]), .A(N1187), .B(N1257));
XOR2XL inst_cellmath__198_0_I834 (.Y(inst_cellmath__198_0_out0[28]), .A(N1189), .B(N1269));
XOR2XL inst_cellmath__198_0_I835 (.Y(inst_cellmath__198_0_out0[32]), .A(N1191), .B(N1281));
XNOR2X1 node_cs_reduced_local_A_I900 (.Y(N1292), .A(N1230), .B(N1034));
XNOR2X1 node_cs_reduced_local_A_I901 (.Y(N1293), .A(N1230), .B(N1033));
MXI2XL inst_cellmath__198_0_I837 (.Y(inst_cellmath__198_0_out0[15]), .A(N1292), .B(N1293), .S0(N1777));
XNOR2X1 node_cs_reduced_local_A_I902 (.Y(N1295), .A(N1236), .B(N1038));
XNOR2X1 node_cs_reduced_local_A_I903 (.Y(N1296), .A(N1236), .B(N1037));
MXI2XL inst_cellmath__198_0_I839 (.Y(inst_cellmath__198_0_out0[17]), .A(N1295), .B(N1296), .S0(N1778));
XNOR2X1 node_cs_reduced_local_A_I904 (.Y(N1298), .A(N1242), .B(N1042));
XNOR2X1 node_cs_reduced_local_A_I1197 (.Y(N1299), .A(N1041), .B(N1242));
MXI2X1 inst_cellmath__198_0_I841 (.Y(inst_cellmath__198_0_out0[19]), .A(N1298), .B(N1299), .S0(N1165));
XNOR2X1 node_cs_reduced_local_A_I906 (.Y(N1301), .A(N1248), .B(N1046));
XNOR2X1 node_cs_reduced_local_A_I907 (.Y(N1302), .A(N1248), .B(N1045));
MXI2XL inst_cellmath__198_0_I843 (.Y(inst_cellmath__198_0_out0[21]), .A(N1301), .B(N1302), .S0(N1167));
XNOR2X1 node_cs_reduced_local_A_I908 (.Y(N1304), .A(N1254), .B(N1050));
XNOR2X1 node_cs_reduced_local_A_I909 (.Y(N1305), .A(N1254), .B(N1049));
MXI2X1 inst_cellmath__198_0_I845 (.Y(inst_cellmath__198_0_out0[23]), .A(N1305), .B(N1304), .S0(N1185));
XNOR2X1 node_cs_reduced_local_A_I910 (.Y(N1307), .A(N1260), .B(N1054));
XNOR2X1 node_cs_reduced_local_A_I911 (.Y(N1308), .A(N1260), .B(N1053));
MXI2XL inst_cellmath__198_0_I847 (.Y(inst_cellmath__198_0_out0[25]), .A(N1308), .B(N1307), .S0(N1187));
XNOR2X1 node_cs_local_A_I912 (.Y(N1310), .A(N1263), .B(N1795));
NOR2BX1 node_cs_local_A_I1198 (.Y(N1529), .AN(N1098), .B(N1795));
XOR2XL node_cs_local_A_I914 (.Y(N1311), .A(N1263), .B(N1529));
MXI2XL inst_cellmath__198_0_I849 (.Y(inst_cellmath__198_0_out0[26]), .A(N1310), .B(N1311), .S0(N1187));
XNOR2X1 node_cs_local_A_I915 (.Y(N1313), .A(N1266), .B(N1107));
NOR2XL node_cs_local_A_I916 (.Y(N1538), .A(N1108), .B(N1107));
XOR2XL node_cs_local_A_I917 (.Y(N1314), .A(N1266), .B(N1538));
MXI2XL inst_cellmath__198_0_I851 (.Y(inst_cellmath__198_0_out0[27]), .A(N1313), .B(N1314), .S0(N1187));
XNOR2X1 node_cs_reduced_local_A_I918 (.Y(N1316), .A(N1272), .B(N1062));
XNOR2X1 node_cs_reduced_local_A_I919 (.Y(N1317), .A(N1272), .B(N1061));
MXI2XL inst_cellmath__198_0_I853 (.Y(inst_cellmath__198_0_out0[29]), .A(N1317), .B(N1316), .S0(N1189));
XNOR2X1 node_cs_local_A_I920 (.Y(N1319), .A(N1275), .B(N1801));
NOR2BX1 node_cs_local_A_I1199 (.Y(N1554), .AN(N1114), .B(N1801));
XOR2XL node_cs_local_A_I922 (.Y(N1320), .A(N1275), .B(N1554));
MXI2XL inst_cellmath__198_0_I855 (.Y(inst_cellmath__198_0_out0[30]), .A(N1319), .B(N1320), .S0(N1189));
XNOR2X1 node_cs_local_A_I923 (.Y(N1322), .A(N1278), .B(N1123));
NOR2XL node_cs_local_A_I924 (.Y(N1563), .A(N1124), .B(N1123));
XOR2XL node_cs_local_A_I925 (.Y(N1323), .A(N1278), .B(N1563));
MXI2XL inst_cellmath__198_0_I857 (.Y(inst_cellmath__198_0_out0[31]), .A(N1322), .B(N1323), .S0(N1189));
assign inst_cellmath__198_0_out0[1] = 1'B0;
endmodule

module cynw_cm_float_sin_inst_cellmath__203_0_bdw1946085813_bdw (
	inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1,
	inst_cellmath__203_0_in0,
	inst_cellmath__203_0_in1,
	inst_cellmath__203_0_in2,
	inst_cellmath__203_0_in3,
	inst_cellmath__203_0_in4
	); /* architecture "gate_level" */ 
output [46:0] inst_cellmath__203_0_out0,
	inst_cellmath__203_0_out1;
input [15:0] inst_cellmath__203_0_in0;
input [32:17] inst_cellmath__203_0_in1;
input [42:23] inst_cellmath__203_0_in2;
input [21:0] inst_cellmath__203_0_in3;
input [0:0] inst_cellmath__203_0_in4;
wire N518,N520,N522,N524,N526,N528,N530 
	,N532,N534,N536,N538,N540,N542,N544,N546 
	,N548,N550,N552,N554,N560,N567,N568,N569 
	,N570,N571,N572,N573,N574,N575,N576,N577 
	,N578,N579,N580,N581,N582,N583,N584,N585 
	,N589,N590,N591,N595,N596,N597,N598,N599 
	,N600,N601,N602,N603,N604,N605,N606,N607 
	,N608,N609,N610,N611,N612,N613,N614,N615 
	,N621,N625,N626,N627,N628,N629,N630,N631 
	,N632,N633,N634,N635,N636,N637,N638,N639 
	,N640,N641,N642,N643,N644,N645,N649,N651 
	,N655,N656,N657,N658,N659,N660,N661,N662 
	,N663,N664,N665,N666,N667,N668,N669,N670 
	,N671,N672,N673,N674,N675,N680,N681,N685 
	,N686,N687,N688,N689,N690,N691,N692,N693 
	,N694,N695,N696,N697,N698,N699,N700,N701 
	,N702,N703,N704,N705,N709,N710,N711,N715 
	,N716,N717,N718,N719,N720,N721,N722,N723 
	,N724,N725,N726,N727,N728,N729,N730,N731 
	,N732,N733,N734,N735,N741,N745,N746,N747 
	,N748,N749,N750,N751,N752,N753,N754,N755 
	,N756,N757,N758,N759,N760,N761,N762,N763 
	,N764,N765,N768,N770,N779,N781,N783,N785 
	,N787,N789,N791,N793,N795,N797,N799,N801 
	,N803,N805,N807,N809,N811,N813,N815,N817 
	,N819,N1025,N1027,N1029,N1031,N1033,N1035,N1037 
	,N1039,N1041,N1043,N1045,N1047,N1049,N1051,N1053 
	,N1055,N1061,N1067,N1077,N1078,N1079,N1080,N1081 
	,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089 
	,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097 
	,N1098,N1099,N1103,N1105,N1109,N1110,N1111,N1112 
	,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120 
	,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128 
	,N1129,N1130,N1131,N1135,N1137,N1141,N1142,N1143 
	,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151 
	,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159 
	,N1160,N1161,N1162,N1163,N1167,N1169,N1173,N1174 
	,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182 
	,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190 
	,N1191,N1192,N1193,N1194,N1195,N1199,N1201,N1205 
	,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213 
	,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221 
	,N1222,N1223,N1224,N1225,N1226,N1227,N1231,N1233 
	,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244 
	,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252 
	,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1263 
	,N1265,N1269,N1270,N1271,N1272,N1273,N1274,N1275 
	,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283 
	,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1295 
	,N1297,N1301,N1302,N1303,N1304,N1305,N1306,N1307 
	,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315 
	,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1366 
	,N1376,N1379,N1380,N1382,N1384,N1387,N1388,N1389 
	,N1390,N1391,N1392,N1395,N1396,N1397,N1398,N1399 
	,N1400,N1403,N1404,N1405,N1406,N1407,N1408,N1409 
	,N1410,N1411,N1412,N1415,N1416,N1417,N1418,N1419 
	,N1420,N1421,N1422,N1423,N1424,N1427,N1428,N1429 
	,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437 
	,N1438,N1439,N1440,N1443,N1444,N1445,N1446,N1447 
	,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455 
	,N1456,N1459,N1460,N1461,N1462,N1463,N1464,N1465 
	,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473 
	,N1474,N1475,N1476,N1479,N1480,N1481,N1482,N1483 
	,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491 
	,N1492,N1493,N1494,N1495,N1496,N1499,N1500,N1501 
	,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509 
	,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517 
	,N1518,N1519,N1520,N1523,N1524,N1525,N1526,N1527 
	,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535 
	,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543 
	,N1544,N1547,N1548,N1549,N1550,N1551,N1552,N1553 
	,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561 
	,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569 
	,N1570,N1571,N1572,N1575,N1576,N1577,N1578,N1579 
	,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587 
	,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595 
	,N1596,N1597,N1598,N1599,N1600,N1603,N1604,N1605 
	,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613 
	,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621 
	,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629 
	,N1630,N1633,N1634,N1635,N1636,N1637,N1638,N1639 
	,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647 
	,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655 
	,N1656,N1657,N1658,N1659,N1660,N1663,N1664,N1665 
	,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673 
	,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681 
	,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689 
	,N1690,N1691,N1692,N1695,N1696,N1698,N1699,N1700 
	,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708 
	,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716 
	,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724 
	,N1725,N1726,N1729,N1730,N1732,N1733,N1734,N1735 
	,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743 
	,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751 
	,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759 
	,N1760,N1763,N1764,N1765,N1766,N1767,N1768,N1769 
	,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777 
	,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785 
	,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1795 
	,N1796,N1798,N1799,N1800,N1801,N1802,N1803,N1804 
	,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812 
	,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820 
	,N1821,N1822,N1823,N1824,N1827,N1828,N1830,N1831 
	,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839 
	,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847 
	,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855 
	,N1856,N1859,N1860,N1863,N1864,N1865,N1866,N1867 
	,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875 
	,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883 
	,N1884,N1885,N1886,N1887,N1888,N1891,N1892,N1893 
	,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901 
	,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909 
	,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1919 
	,N1920,N1923,N1924,N1925,N1926,N1927,N1928,N1929 
	,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937 
	,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1947 
	,N1948,N1951,N1952,N1953,N1954,N1955,N1956,N1957 
	,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965 
	,N1966,N1967,N1968,N1969,N1970,N1973,N1974,N1975 
	,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983 
	,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991 
	,N1992,N1995,N1996,N1999,N2000,N2001,N2002,N2003 
	,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011 
	,N2012,N2013,N2014,N2017,N2018,N2019,N2020,N2021 
	,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029 
	,N2030,N2031,N2032,N2035,N2036,N2039,N2040,N2041 
	,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049 
	,N2050,N2053,N2054,N2055,N2056,N2057,N2058,N2059 
	,N2060,N2061,N2062,N2063,N2064,N2067,N2068,N2071 
	,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2081 
	,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2091 
	,N2092,N2095,N2096,N2097,N2098,N2101,N2102,N2103 
	,N2104,N2107,N2108,N2111,N2112,N2226,N2235,N2244 
	,N2253,N2262,N2271,N2280,N2289,N2298,N2307,N2316 
	,N2325,N2334,N2343,N2352,N2361,N2370,N2379,N2388 
	,N2397,N2406,N2415,N2417,N2428,N2437,N2446,N2455 
	,N2464,N2473,N2482,N2491,N2500,N2509,N2518,N2527 
	,N2536,N2545,N2554,N2563,N2572,N2581,N2590,N2599 
	,N2608,N2617,N2619,N2630,N2639,N2648,N2657,N2666 
	,N2675,N2684,N2693,N2702,N2711,N2720,N2729,N2738 
	,N2747,N2756,N2765,N2774,N2783,N2792,N2801,N2810 
	,N2819,N2821,N2832,N2841,N2850,N2859,N2868,N2877 
	,N2886,N2895,N2904,N2913,N2922,N2931,N2940,N2949 
	,N2958,N2967,N2976,N2985,N2994,N3003,N3012,N3021 
	,N3023,N3034,N3043,N3052,N3061,N3070,N3079,N3088 
	,N3097,N3106,N3115,N3124,N3133,N3142,N3151,N3160 
	,N3169,N3178,N3187,N3196,N3205,N3214,N3223,N3225 
	,N3236,N3245,N3254,N3263,N3272,N3281,N3290,N3299 
	,N3308,N3317,N3326,N3335,N3344,N3353,N3362,N3371 
	,N3380,N3389,N3398,N3407,N3416,N3425,N3427,N3438 
	,N3447,N3456,N3465,N3474,N3483,N3492,N3501,N3510 
	,N3519,N3528,N3537,N3546,N3555,N3564,N3573,N3582 
	,N3591,N3600,N3609,N3618,N3640,N3649,N3658,N3667 
	,N3676,N3685,N3694,N3703,N3712,N3721,N3730,N3739 
	,N3748,N3757,N3766,N3775,N3784,N3793,N3802,N3811 
	,N3820,N3829,N3838,N3847,N3849,N3860,N3869,N3878 
	,N3887,N3896,N3905,N3914,N3923,N3932,N3941,N3950 
	,N3959,N3968,N3977,N3986,N3995,N4004,N4013,N4022 
	,N4031,N4040,N4049,N4058,N4067,N4069,N4080,N4089 
	,N4098,N4107,N4116,N4125,N4134,N4143,N4152,N4161 
	,N4170,N4179,N4188,N4197,N4206,N4215,N4224,N4233 
	,N4242,N4251,N4260,N4269,N4278,N4287,N4289,N4300 
	,N4309,N4318,N4327,N4336,N4345,N4354,N4363,N4372 
	,N4381,N4390,N4399,N4408,N4417,N4426,N4435,N4444 
	,N4453,N4462,N4471,N4480,N4489,N4498,N4507,N4509 
	,N4520,N4529,N4538,N4547,N4556,N4565,N4574,N4583 
	,N4592,N4601,N4610,N4619,N4628,N4637,N4646,N4655 
	,N4664,N4673,N4682,N4691,N4700,N4709,N4718,N4727 
	,N4729,N4740,N4749,N4758,N4767,N4776,N4785,N4794 
	,N4803,N4812,N4821,N4830,N4839,N4848,N4857,N4866 
	,N4875,N4884,N4893,N4902,N4911,N4920,N4929,N4938 
	,N4947,N4949,N4960,N4969,N4978,N4987,N4996,N5005 
	,N5014,N5023,N5032,N5041,N5050,N5059,N5068,N5077 
	,N5086,N5095,N5104,N5113,N5122,N5131,N5140,N5149 
	,N5158,N5167,N5169,N5180,N5189,N5198,N5207,N5216 
	,N5225,N5234,N5243,N5252,N5261,N5270,N5279,N5288 
	,N5297,N5306,N5315,N5324,N5333,N5342,N5351,N5360 
	,N5369,N5378,N5387,N5396,N5405,N5414,N5435,N5444 
	,N5453,N5462,N5471,N5617,N5624,N5625,N5626,N5627 
	,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635 
	,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5644 
	,N5645,N5647,N5649,N5650,N5654,N5658,N5666,N5667 
	,N5668,N5670,N5671,N5672,N5673,N5674,N5675,N5681 
	,N5683,N5684,N5685,N5686,N5687,N5688,N5689,N5698 
	,N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5713 
	,N5719,N5721,N5722,N5723,N5729,N5731,N5732,N5733 
	,N5736,N5737,N5738,N5739,N5745,N5747,N5748,N5749 
	,N5754,N5755,N5763,N5764,N5765,N5766,N5767,N5768 
	,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776 
	,N5777,N5778,N5779,N5780,N5781,N5782,N5783,N5784 
	,N5785,N5786,N5787,N5788,N5789,N5797,N5805,N5806 
	,N5815,N5816,N5817,N5818,N5833,N5842,N5843,N5844 
	,N5859,N5868,N5869,N5870,N5871,N5872,N5887,N5896 
	,N5897,N5898,N5899,N5900,N5915,N5924,N5939,N5947 
	,N5962,N5970,N5985;
INVXL inst_cellmath__203_0_I1819 (.Y(N5617), .A(inst_cellmath__203_0_in2[23]));
INVXL inst_cellmath__203_0_I1826 (.Y(N5624), .A(inst_cellmath__203_0_in2[24]));
INVXL inst_cellmath__203_0_I1827 (.Y(N5625), .A(inst_cellmath__203_0_in2[25]));
INVXL inst_cellmath__203_0_I1828 (.Y(N5626), .A(inst_cellmath__203_0_in2[26]));
INVXL inst_cellmath__203_0_I1829 (.Y(N5627), .A(inst_cellmath__203_0_in2[27]));
INVXL inst_cellmath__203_0_I1830 (.Y(N5628), .A(inst_cellmath__203_0_in2[28]));
INVXL inst_cellmath__203_0_I1831 (.Y(N5629), .A(inst_cellmath__203_0_in2[29]));
INVXL inst_cellmath__203_0_I1832 (.Y(N5630), .A(inst_cellmath__203_0_in2[30]));
INVXL inst_cellmath__203_0_I1833 (.Y(N5631), .A(inst_cellmath__203_0_in2[31]));
INVXL inst_cellmath__203_0_I1834 (.Y(N5632), .A(inst_cellmath__203_0_in2[32]));
INVXL inst_cellmath__203_0_I1835 (.Y(N5633), .A(inst_cellmath__203_0_in2[33]));
INVXL inst_cellmath__203_0_I1836 (.Y(N5634), .A(inst_cellmath__203_0_in2[34]));
INVXL inst_cellmath__203_0_I1837 (.Y(N5635), .A(inst_cellmath__203_0_in2[35]));
INVXL inst_cellmath__203_0_I1838 (.Y(N5636), .A(inst_cellmath__203_0_in2[36]));
INVXL inst_cellmath__203_0_I1839 (.Y(N5637), .A(inst_cellmath__203_0_in2[37]));
INVXL inst_cellmath__203_0_I1840 (.Y(N5638), .A(inst_cellmath__203_0_in2[38]));
INVXL inst_cellmath__203_0_I1841 (.Y(N5639), .A(inst_cellmath__203_0_in2[39]));
INVXL inst_cellmath__203_0_I1842 (.Y(N5640), .A(inst_cellmath__203_0_in2[40]));
INVXL inst_cellmath__203_0_I1843 (.Y(N5641), .A(inst_cellmath__203_0_in2[41]));
INVXL inst_cellmath__203_0_I1844 (.Y(N5642), .A(inst_cellmath__203_0_in2[42]));
BUFX6 inst_cellmath__203_0_I2205 (.Y(N5644), .A(inst_cellmath__203_0_in1[17]));
INVXL inst_cellmath__203_0_I1852 (.Y(N5650), .A(N5644));
INVXL inst_cellmath__203_0_I1851 (.Y(N5649), .A(N5644));
INVXL inst_cellmath__203_0_I1849 (.Y(N5647), .A(N5644));
INVX2 inst_cellmath__203_0_I1847 (.Y(N5645), .A(N5644));
NOR2XL inst_cellmath__203_0_I71 (.Y(inst_cellmath__203_0_out1[0]), .A(N5649), .B(N5617));
NOR2XL inst_cellmath__203_0_I72 (.Y(N518), .A(N5649), .B(N5624));
NOR2XL inst_cellmath__203_0_I73 (.Y(N520), .A(N5649), .B(N5625));
NOR2XL inst_cellmath__203_0_I74 (.Y(N522), .A(N5649), .B(N5626));
NOR2XL inst_cellmath__203_0_I75 (.Y(N524), .A(N5649), .B(N5627));
NOR2XL inst_cellmath__203_0_I76 (.Y(N526), .A(N5649), .B(N5628));
NOR2XL inst_cellmath__203_0_I77 (.Y(N528), .A(N5649), .B(N5629));
NOR2XL inst_cellmath__203_0_I78 (.Y(N530), .A(N5649), .B(N5630));
NOR2XL inst_cellmath__203_0_I79 (.Y(N532), .A(N5647), .B(N5631));
NOR2XL inst_cellmath__203_0_I80 (.Y(N534), .A(N5647), .B(N5632));
NOR2XL inst_cellmath__203_0_I81 (.Y(N536), .A(N5647), .B(N5633));
NOR2XL inst_cellmath__203_0_I82 (.Y(N538), .A(N5647), .B(N5634));
NOR2XL inst_cellmath__203_0_I83 (.Y(N540), .A(N5650), .B(N5635));
NOR2XL inst_cellmath__203_0_I84 (.Y(N542), .A(N5650), .B(N5636));
NOR2XL inst_cellmath__203_0_I85 (.Y(N544), .A(N5650), .B(N5637));
NOR2XL inst_cellmath__203_0_I86 (.Y(N546), .A(N5650), .B(N5638));
NOR2XL inst_cellmath__203_0_I87 (.Y(N548), .A(N5645), .B(N5639));
NOR2XL inst_cellmath__203_0_I88 (.Y(N550), .A(N5645), .B(N5640));
NOR2XL inst_cellmath__203_0_I89 (.Y(N552), .A(N5645), .B(N5641));
NOR2XL inst_cellmath__203_0_I90 (.Y(N554), .A(N5645), .B(N5642));
NOR2BX1 inst_cellmath__203_0_I1817 (.Y(N560), .AN(inst_cellmath__203_0_in1[18]), .B(inst_cellmath__203_0_in1[19]));
INVXL inst_cellmath__203_0_I1860 (.Y(N5658), .A(inst_cellmath__203_0_in1[18]));
INVXL inst_cellmath__203_0_I1856 (.Y(N5654), .A(inst_cellmath__203_0_in1[18]));
INVX1 inst_cellmath__203_0_I1868 (.Y(N5666), .A(N560));
INVXL inst_cellmath__203_0_I1869 (.Y(N5667), .A(inst_cellmath__203_0_in1[19]));
NOR2XL addgen2_A_I1059 (.Y(N2226), .A(N5617), .B(N5654));
MXI2X2 addgen2_A_I1060 (.Y(inst_cellmath__203_0_out1[1]), .A(N5667), .B(N5666), .S0(N2226));
MXI2XL inst_cellmath__203_0_I1061 (.Y(N2235), .A(N5624), .B(N5617), .S0(N5658));
MX2XL inst_cellmath__203_0_I2207 (.Y(N5668), .A(N5667), .B(N5666), .S0(N2235));
INVXL inst_cellmath__203_0_I1871 (.Y(inst_cellmath__203_0_out1[2]), .A(N5668));
MXI2XL addgen2_A_I1063 (.Y(N2244), .A(N5625), .B(N5624), .S0(N5658));
MXI2XL addgen2_A_I1064 (.Y(N567), .A(N5667), .B(N5666), .S0(N2244));
MXI2XL addgen2_A_I1065 (.Y(N2253), .A(N5626), .B(N5625), .S0(N5658));
MXI2XL addgen2_A_I1066 (.Y(N568), .A(N5667), .B(N5666), .S0(N2253));
MXI2XL addgen2_A_I1067 (.Y(N2262), .A(N5627), .B(N5626), .S0(N5658));
MXI2XL addgen2_A_I1068 (.Y(N569), .A(N5667), .B(N5666), .S0(N2262));
MXI2XL addgen2_A_I1069 (.Y(N2271), .A(N5628), .B(N5627), .S0(N5658));
MXI2XL addgen2_A_I1070 (.Y(N570), .A(N5667), .B(N5666), .S0(N2271));
MXI2XL addgen2_A_I1071 (.Y(N2280), .A(N5629), .B(N5628), .S0(N5658));
MXI2XL addgen2_A_I1072 (.Y(N571), .A(N5667), .B(N5666), .S0(N2280));
MXI2XL addgen2_A_I1073 (.Y(N2289), .A(N5630), .B(N5629), .S0(N5658));
MXI2XL addgen2_A_I1074 (.Y(N572), .A(N5667), .B(N5666), .S0(N2289));
MXI2XL addgen2_A_I1075 (.Y(N2298), .A(N5631), .B(N5630), .S0(N5658));
MXI2XL addgen2_A_I1076 (.Y(N573), .A(N5667), .B(N5666), .S0(N2298));
MXI2XL addgen2_A_I1077 (.Y(N2307), .A(N5632), .B(N5631), .S0(N5658));
MXI2XL addgen2_A_I1078 (.Y(N574), .A(N5667), .B(N5666), .S0(N2307));
MXI2XL addgen2_A_I1079 (.Y(N2316), .A(N5633), .B(N5632), .S0(N5658));
MXI2XL addgen2_A_I1080 (.Y(N575), .A(N5667), .B(N5666), .S0(N2316));
MXI2XL addgen2_A_I1081 (.Y(N2325), .A(N5634), .B(N5633), .S0(N5658));
MXI2XL addgen2_A_I1082 (.Y(N576), .A(N5667), .B(N5666), .S0(N2325));
MXI2XL addgen2_A_I1083 (.Y(N2334), .A(N5635), .B(N5634), .S0(N5658));
MXI2XL addgen2_A_I1084 (.Y(N577), .A(N5667), .B(N5666), .S0(N2334));
MXI2XL addgen2_A_I1085 (.Y(N2343), .A(N5636), .B(N5635), .S0(N5658));
MXI2XL addgen2_A_I1086 (.Y(N578), .A(N5667), .B(N5666), .S0(N2343));
MXI2XL addgen2_A_I1087 (.Y(N2352), .A(N5637), .B(N5636), .S0(N5654));
MXI2XL addgen2_A_I1088 (.Y(N579), .A(N5667), .B(N5666), .S0(N2352));
MXI2XL addgen2_A_I1089 (.Y(N2361), .A(N5638), .B(N5637), .S0(N5654));
MXI2XL addgen2_A_I1090 (.Y(N580), .A(N5667), .B(N5666), .S0(N2361));
MXI2XL addgen2_A_I1091 (.Y(N2370), .A(N5639), .B(N5638), .S0(N5654));
MXI2XL addgen2_A_I1092 (.Y(N581), .A(N5667), .B(N5666), .S0(N2370));
MXI2XL addgen2_A_I1093 (.Y(N2379), .A(N5640), .B(N5639), .S0(N5654));
MXI2XL addgen2_A_I1094 (.Y(N582), .A(N5667), .B(N5666), .S0(N2379));
MXI2XL addgen2_A_I1095 (.Y(N2388), .A(N5641), .B(N5640), .S0(N5654));
MXI2XL addgen2_A_I1096 (.Y(N583), .A(N5667), .B(N5666), .S0(N2388));
MXI2XL addgen2_A_I1097 (.Y(N2397), .A(N5642), .B(N5641), .S0(N5654));
MXI2XL addgen2_A_I1098 (.Y(N584), .A(N5667), .B(N5666), .S0(N2397));
NAND2XL addgen2_A_I1099 (.Y(N2406), .A(N5642), .B(N5654));
MXI2XL addgen2_A_I1100 (.Y(N585), .A(N5667), .B(N5666), .S0(N2406));
XNOR2X1 enc2_A_I1101 (.Y(N589), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
NAND2XL enc2_A_I1102 (.Y(N2415), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
NOR2XL enc2_A_I1103 (.Y(N2417), .A(inst_cellmath__203_0_in1[20]), .B(inst_cellmath__203_0_in1[19]));
AND2XL enc2_A_I1104 (.Y(N591), .A(N2415), .B(inst_cellmath__203_0_in1[21]));
NOR2XL enc2_A_I1105 (.Y(N590), .A(N2417), .B(inst_cellmath__203_0_in1[21]));
INVX3 inst_cellmath__203_0_I1872 (.Y(N5670), .A(N589));
INVXL inst_cellmath__203_0_I1877 (.Y(N5675), .A(N5670));
INVX2 inst_cellmath__203_0_I1876 (.Y(N5674), .A(N5670));
INVX1 inst_cellmath__203_0_I1875 (.Y(N5673), .A(N5670));
INVX1 inst_cellmath__203_0_I1874 (.Y(N5672), .A(N5670));
INVX2 inst_cellmath__203_0_I1873 (.Y(N5671), .A(N5670));
INVX2 inst_cellmath__203_0_I1885 (.Y(N5683), .A(N590));
INVXL inst_cellmath__203_0_I1883 (.Y(N5681), .A(N590));
INVX2 inst_cellmath__203_0_I1886 (.Y(N5684), .A(N591));
NOR2XL addgen2_A_I1106 (.Y(N2428), .A(N5617), .B(N5671));
MXI2XL addgen2_A_I1107 (.Y(N595), .A(N5684), .B(N5683), .S0(N2428));
MXI2XL addgen2_A_I1108 (.Y(N2437), .A(N5624), .B(N5617), .S0(N5675));
MXI2XL addgen2_A_I1109 (.Y(N596), .A(N5684), .B(N5683), .S0(N2437));
MXI2X1 addgen2_A_I1110 (.Y(N2446), .A(N5625), .B(N5624), .S0(N5674));
MXI2X1 addgen2_A_I1111 (.Y(N597), .A(N5684), .B(N5683), .S0(N2446));
MXI2XL addgen2_A_I1112 (.Y(N2455), .A(N5626), .B(N5625), .S0(N5674));
MXI2XL addgen2_A_I1113 (.Y(N598), .A(N5684), .B(N5683), .S0(N2455));
MXI2XL addgen2_A_I1114 (.Y(N2464), .A(N5627), .B(N5626), .S0(N5674));
MXI2XL addgen2_A_I1115 (.Y(N599), .A(N5684), .B(N5683), .S0(N2464));
MXI2XL addgen2_A_I1116 (.Y(N2473), .A(N5628), .B(N5627), .S0(N5674));
MXI2XL addgen2_A_I1117 (.Y(N600), .A(N5684), .B(N5681), .S0(N2473));
MXI2XL addgen2_A_I1118 (.Y(N2482), .A(N5629), .B(N5628), .S0(N5674));
MXI2XL addgen2_A_I1119 (.Y(N601), .A(N5684), .B(N5681), .S0(N2482));
MXI2XL addgen2_A_I1120 (.Y(N2491), .A(N5630), .B(N5629), .S0(N5673));
MXI2XL addgen2_A_I1121 (.Y(N602), .A(N5684), .B(N5681), .S0(N2491));
MXI2XL addgen2_A_I1122 (.Y(N2500), .A(N5631), .B(N5630), .S0(N5673));
MXI2XL addgen2_A_I1123 (.Y(N603), .A(N5684), .B(N5681), .S0(N2500));
MXI2XL addgen2_A_I1124 (.Y(N2509), .A(N5632), .B(N5631), .S0(N5673));
MXI2XL addgen2_A_I1125 (.Y(N604), .A(N5684), .B(N5681), .S0(N2509));
MXI2XL addgen2_A_I1126 (.Y(N2518), .A(N5633), .B(N5632), .S0(N5673));
MXI2XL addgen2_A_I1127 (.Y(N605), .A(N5684), .B(N5681), .S0(N2518));
MXI2X1 addgen2_A_I1128 (.Y(N2527), .A(N5634), .B(N5633), .S0(N5673));
MXI2X1 addgen2_A_I1129 (.Y(N606), .A(N5684), .B(N5681), .S0(N2527));
MXI2XL addgen2_A_I1130 (.Y(N2536), .A(N5635), .B(N5634), .S0(N5672));
MXI2XL addgen2_A_I1131 (.Y(N607), .A(N5684), .B(N5681), .S0(N2536));
MXI2XL addgen2_A_I1132 (.Y(N2545), .A(N5636), .B(N5635), .S0(N5672));
MXI2XL addgen2_A_I1133 (.Y(N608), .A(N5684), .B(N5683), .S0(N2545));
MXI2XL addgen2_A_I1134 (.Y(N2554), .A(N5637), .B(N5636), .S0(N5672));
MXI2XL addgen2_A_I1135 (.Y(N609), .A(N5684), .B(N5683), .S0(N2554));
MXI2XL addgen2_A_I1136 (.Y(N2563), .A(N5638), .B(N5637), .S0(N5672));
MXI2XL addgen2_A_I1137 (.Y(N610), .A(N5684), .B(N5683), .S0(N2563));
MXI2X1 addgen2_A_I1138 (.Y(N2572), .A(N5639), .B(N5638), .S0(N5672));
MXI2X1 addgen2_A_I1139 (.Y(N611), .A(N5684), .B(N5683), .S0(N2572));
MXI2XL addgen2_A_I1140 (.Y(N2581), .A(N5640), .B(N5639), .S0(N5671));
MXI2XL addgen2_A_I1141 (.Y(N612), .A(N5684), .B(N5683), .S0(N2581));
MXI2XL addgen2_A_I1142 (.Y(N2590), .A(N5641), .B(N5640), .S0(N5671));
MXI2XL addgen2_A_I1143 (.Y(N613), .A(N5684), .B(N5683), .S0(N2590));
MXI2X1 addgen2_A_I1144 (.Y(N2599), .A(N5642), .B(N5641), .S0(N5671));
MXI2X1 addgen2_A_I1145 (.Y(N614), .A(N5684), .B(N5683), .S0(N2599));
NAND2XL addgen2_A_I1146 (.Y(N2608), .A(N5642), .B(N5671));
MXI2XL addgen2_A_I1147 (.Y(N615), .A(N5684), .B(N5683), .S0(N2608));
NAND2XL enc2_A_I1149 (.Y(N2617), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
NOR2XL enc2_A_I1150 (.Y(N2619), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
AND2XL enc2_A_I1151 (.Y(N621), .A(N2617), .B(inst_cellmath__203_0_in1[23]));
CLKXOR2X1 inst_cellmath__203_0_I2200 (.Y(N5685), .A(inst_cellmath__203_0_in1[22]), .B(inst_cellmath__203_0_in1[21]));
INVXL inst_cellmath__203_0_I1891 (.Y(N5689), .A(N5685));
INVX1 inst_cellmath__203_0_I1890 (.Y(N5688), .A(N5685));
INVX1 inst_cellmath__203_0_I1889 (.Y(N5687), .A(N5685));
INVX1 inst_cellmath__203_0_I1888 (.Y(N5686), .A(N5685));
OR2X2 inst_cellmath__203_0_I2211 (.Y(N5698), .A(N2619), .B(inst_cellmath__203_0_in1[23]));
INVX2 inst_cellmath__203_0_I1901 (.Y(N5699), .A(N621));
NOR2X1 addgen2_A_I1153 (.Y(N2630), .A(N5617), .B(N5686));
MXI2X1 addgen2_A_I1154 (.Y(N625), .A(N5699), .B(N5698), .S0(N2630));
MXI2XL addgen2_A_I2212 (.Y(N2639), .A(N5617), .B(N5624), .S0(N5685));
MXI2XL addgen2_A_I1156 (.Y(N626), .A(N5699), .B(N5698), .S0(N2639));
MXI2XL addgen2_A_I1157 (.Y(N2648), .A(N5625), .B(N5624), .S0(N5689));
MXI2XL addgen2_A_I1158 (.Y(N627), .A(N5699), .B(N5698), .S0(N2648));
MXI2XL addgen2_A_I1159 (.Y(N2657), .A(N5626), .B(N5625), .S0(N5689));
MXI2XL addgen2_A_I1160 (.Y(N628), .A(N5699), .B(N5698), .S0(N2657));
MXI2XL addgen2_A_I1161 (.Y(N2666), .A(N5627), .B(N5626), .S0(N5689));
MXI2XL addgen2_A_I1162 (.Y(N629), .A(N5699), .B(N5698), .S0(N2666));
MXI2XL addgen2_A_I1163 (.Y(N2675), .A(N5628), .B(N5627), .S0(N5689));
MXI2XL addgen2_A_I1164 (.Y(N630), .A(N5699), .B(N5698), .S0(N2675));
MXI2XL addgen2_A_I1165 (.Y(N2684), .A(N5629), .B(N5628), .S0(N5689));
MXI2XL addgen2_A_I1166 (.Y(N631), .A(N5699), .B(N5698), .S0(N2684));
MXI2XL addgen2_A_I1167 (.Y(N2693), .A(N5630), .B(N5629), .S0(N5688));
MXI2XL addgen2_A_I1168 (.Y(N632), .A(N5699), .B(N5698), .S0(N2693));
MXI2XL addgen2_A_I1169 (.Y(N2702), .A(N5631), .B(N5630), .S0(N5688));
MXI2XL addgen2_A_I1170 (.Y(N633), .A(N5699), .B(N5698), .S0(N2702));
MXI2XL addgen2_A_I1171 (.Y(N2711), .A(N5632), .B(N5631), .S0(N5688));
MXI2XL addgen2_A_I1172 (.Y(N634), .A(N5699), .B(N5698), .S0(N2711));
MXI2XL addgen2_A_I1173 (.Y(N2720), .A(N5633), .B(N5632), .S0(N5688));
MXI2XL addgen2_A_I1174 (.Y(N635), .A(N5699), .B(N5698), .S0(N2720));
MXI2XL addgen2_A_I1175 (.Y(N2729), .A(N5634), .B(N5633), .S0(N5688));
MXI2XL addgen2_A_I1176 (.Y(N636), .A(N5699), .B(N5698), .S0(N2729));
MXI2XL addgen2_A_I1177 (.Y(N2738), .A(N5635), .B(N5634), .S0(N5687));
MXI2XL addgen2_A_I1178 (.Y(N637), .A(N5699), .B(N5698), .S0(N2738));
MXI2XL addgen2_A_I1179 (.Y(N2747), .A(N5636), .B(N5635), .S0(N5687));
MXI2XL addgen2_A_I1180 (.Y(N638), .A(N5699), .B(N5698), .S0(N2747));
MXI2XL addgen2_A_I1181 (.Y(N2756), .A(N5637), .B(N5636), .S0(N5687));
MXI2XL addgen2_A_I1182 (.Y(N639), .A(N5699), .B(N5698), .S0(N2756));
MXI2XL addgen2_A_I1183 (.Y(N2765), .A(N5638), .B(N5637), .S0(N5687));
MXI2XL addgen2_A_I1184 (.Y(N640), .A(N5699), .B(N5698), .S0(N2765));
MXI2XL addgen2_A_I1185 (.Y(N2774), .A(N5639), .B(N5638), .S0(N5687));
MXI2XL addgen2_A_I1186 (.Y(N641), .A(N5699), .B(N5698), .S0(N2774));
MXI2XL addgen2_A_I1187 (.Y(N2783), .A(N5640), .B(N5639), .S0(N5686));
MXI2XL addgen2_A_I1188 (.Y(N642), .A(N5699), .B(N5698), .S0(N2783));
MXI2XL addgen2_A_I1189 (.Y(N2792), .A(N5641), .B(N5640), .S0(N5686));
MXI2XL addgen2_A_I1190 (.Y(N643), .A(N5699), .B(N5698), .S0(N2792));
MXI2XL addgen2_A_I1191 (.Y(N2801), .A(N5642), .B(N5641), .S0(N5686));
MXI2XL addgen2_A_I1192 (.Y(N644), .A(N5699), .B(N5698), .S0(N2801));
NAND2XL addgen2_A_I1193 (.Y(N2810), .A(N5642), .B(N5686));
MXI2XL addgen2_A_I1194 (.Y(N645), .A(N5699), .B(N5698), .S0(N2810));
XNOR2X1 enc2_A_I1195 (.Y(N649), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
NAND2XL enc2_A_I1196 (.Y(N2819), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
NOR2XL enc2_A_I1197 (.Y(N2821), .A(inst_cellmath__203_0_in1[24]), .B(inst_cellmath__203_0_in1[23]));
AND2XL enc2_A_I1198 (.Y(N651), .A(N2819), .B(inst_cellmath__203_0_in1[25]));
INVX3 inst_cellmath__203_0_I1902 (.Y(N5700), .A(N649));
INVXL inst_cellmath__203_0_I1907 (.Y(N5705), .A(N5700));
INVXL inst_cellmath__203_0_I1906 (.Y(N5704), .A(N5700));
INVX2 inst_cellmath__203_0_I1905 (.Y(N5703), .A(N5700));
INVX2 inst_cellmath__203_0_I1904 (.Y(N5702), .A(N5700));
INVXL inst_cellmath__203_0_I1903 (.Y(N5701), .A(N5700));
OR2X1 inst_cellmath__203_0_I2214 (.Y(N5713), .A(N2821), .B(inst_cellmath__203_0_in1[25]));
INVX1 inst_cellmath__203_0_I1923 (.Y(N5721), .A(N651));
INVXL inst_cellmath__203_0_I1921 (.Y(N5719), .A(N651));
NOR2XL addgen2_A_I1200 (.Y(N2832), .A(N5617), .B(N5701));
MXI2XL addgen2_A_I1201 (.Y(N655), .A(N5721), .B(N5713), .S0(N2832));
MXI2XL addgen2_A_I1202 (.Y(N2841), .A(N5624), .B(N5617), .S0(N5705));
MXI2XL addgen2_A_I1203 (.Y(N656), .A(N5721), .B(N5713), .S0(N2841));
MXI2XL addgen2_A_I1204 (.Y(N2850), .A(N5625), .B(N5624), .S0(N5704));
MXI2XL addgen2_A_I1205 (.Y(N657), .A(N5721), .B(N5713), .S0(N2850));
MXI2XL addgen2_A_I1206 (.Y(N2859), .A(N5626), .B(N5625), .S0(N5704));
MXI2XL addgen2_A_I1207 (.Y(N658), .A(N5721), .B(N5713), .S0(N2859));
MXI2XL addgen2_A_I1208 (.Y(N2868), .A(N5627), .B(N5626), .S0(N5704));
MXI2XL addgen2_A_I1209 (.Y(N659), .A(N5721), .B(N5713), .S0(N2868));
MXI2XL addgen2_A_I1210 (.Y(N2877), .A(N5628), .B(N5627), .S0(N5704));
MXI2XL addgen2_A_I1211 (.Y(N660), .A(N5719), .B(N5713), .S0(N2877));
MXI2XL addgen2_A_I1212 (.Y(N2886), .A(N5629), .B(N5628), .S0(N5704));
MXI2XL addgen2_A_I1213 (.Y(N661), .A(N5719), .B(N5713), .S0(N2886));
MXI2XL addgen2_A_I1214 (.Y(N2895), .A(N5630), .B(N5629), .S0(N5703));
MXI2X1 addgen2_A_I1215 (.Y(N662), .A(N5719), .B(N5713), .S0(N2895));
MXI2XL addgen2_A_I1216 (.Y(N2904), .A(N5631), .B(N5630), .S0(N5703));
MXI2XL addgen2_A_I1217 (.Y(N663), .A(N5719), .B(N5713), .S0(N2904));
MXI2XL addgen2_A_I1218 (.Y(N2913), .A(N5632), .B(N5631), .S0(N5703));
MXI2XL addgen2_A_I1219 (.Y(N664), .A(N5721), .B(N5713), .S0(N2913));
MXI2X1 addgen2_A_I1220 (.Y(N2922), .A(N5633), .B(N5632), .S0(N5703));
MXI2X1 addgen2_A_I1221 (.Y(N665), .A(N5721), .B(N5713), .S0(N2922));
MXI2XL addgen2_A_I1222 (.Y(N2931), .A(N5634), .B(N5633), .S0(N5703));
MXI2XL addgen2_A_I1223 (.Y(N666), .A(N5721), .B(N5713), .S0(N2931));
MXI2XL addgen2_A_I1224 (.Y(N2940), .A(N5635), .B(N5634), .S0(N5702));
MXI2XL addgen2_A_I1225 (.Y(N667), .A(N5721), .B(N5713), .S0(N2940));
MXI2XL addgen2_A_I1226 (.Y(N2949), .A(N5636), .B(N5635), .S0(N5702));
MXI2XL addgen2_A_I1227 (.Y(N668), .A(N5721), .B(N5713), .S0(N2949));
MXI2XL addgen2_A_I1228 (.Y(N2958), .A(N5637), .B(N5636), .S0(N5702));
MXI2X1 addgen2_A_I1229 (.Y(N669), .A(N5721), .B(N5713), .S0(N2958));
MXI2X1 addgen2_A_I1230 (.Y(N2967), .A(N5638), .B(N5637), .S0(N5702));
MXI2X1 addgen2_A_I1231 (.Y(N670), .A(N5721), .B(N5713), .S0(N2967));
MXI2XL addgen2_A_I1232 (.Y(N2976), .A(N5639), .B(N5638), .S0(N5702));
MXI2XL addgen2_A_I1233 (.Y(N671), .A(N5721), .B(N5713), .S0(N2976));
MXI2XL addgen2_A_I1234 (.Y(N2985), .A(N5640), .B(N5639), .S0(N5701));
MXI2XL addgen2_A_I1235 (.Y(N672), .A(N5719), .B(N5713), .S0(N2985));
MXI2XL addgen2_A_I1236 (.Y(N2994), .A(N5641), .B(N5640), .S0(N5701));
MXI2XL addgen2_A_I1237 (.Y(N673), .A(N5719), .B(N5713), .S0(N2994));
MXI2XL addgen2_A_I1238 (.Y(N3003), .A(N5642), .B(N5641), .S0(N5701));
MXI2XL addgen2_A_I1239 (.Y(N674), .A(N5719), .B(N5713), .S0(N3003));
NAND2XL addgen2_A_I1240 (.Y(N3012), .A(N5642), .B(N5701));
MXI2XL addgen2_A_I1241 (.Y(N675), .A(N5719), .B(N5713), .S0(N3012));
NAND2XL enc2_A_I1243 (.Y(N3021), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
NOR2XL enc2_A_I1244 (.Y(N3023), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
AND2XL enc2_A_I1245 (.Y(N681), .A(N3021), .B(inst_cellmath__203_0_in1[27]));
NOR2XL enc2_A_I1246 (.Y(N680), .A(N3023), .B(inst_cellmath__203_0_in1[27]));
XOR2XL inst_cellmath__203_0_I2201 (.Y(N5722), .A(inst_cellmath__203_0_in1[26]), .B(inst_cellmath__203_0_in1[25]));
INVX3 inst_cellmath__203_0_I1925 (.Y(N5723), .A(N5722));
INVXL inst_cellmath__203_0_I1933 (.Y(N5731), .A(N680));
INVXL inst_cellmath__203_0_I1931 (.Y(N5729), .A(N680));
INVX2 inst_cellmath__203_0_I1934 (.Y(N5732), .A(N681));
NOR2XL addgen2_A_I1247 (.Y(N3034), .A(N5617), .B(N5723));
MXI2XL addgen2_A_I1248 (.Y(N685), .A(N5732), .B(N5731), .S0(N3034));
MXI2XL addgen2_A_I1249 (.Y(N3043), .A(N5624), .B(N5617), .S0(N5723));
MXI2XL addgen2_A_I1250 (.Y(N686), .A(N5732), .B(N5731), .S0(N3043));
MXI2XL addgen2_A_I1251 (.Y(N3052), .A(N5625), .B(N5624), .S0(N5723));
MXI2XL addgen2_A_I1252 (.Y(N687), .A(N5732), .B(N5731), .S0(N3052));
MXI2XL addgen2_A_I1253 (.Y(N3061), .A(N5626), .B(N5625), .S0(N5723));
MXI2XL addgen2_A_I1254 (.Y(N688), .A(N5732), .B(N5731), .S0(N3061));
MXI2XL addgen2_A_I1255 (.Y(N3070), .A(N5627), .B(N5626), .S0(N5723));
MXI2XL addgen2_A_I1256 (.Y(N689), .A(N5732), .B(N5731), .S0(N3070));
MXI2XL addgen2_A_I1257 (.Y(N3079), .A(N5628), .B(N5627), .S0(N5723));
MXI2XL addgen2_A_I1258 (.Y(N690), .A(N5732), .B(N5729), .S0(N3079));
MXI2XL addgen2_A_I1259 (.Y(N3088), .A(N5629), .B(N5628), .S0(N5723));
MXI2XL addgen2_A_I1260 (.Y(N691), .A(N5732), .B(N5729), .S0(N3088));
MXI2XL addgen2_A_I1261 (.Y(N3097), .A(N5630), .B(N5629), .S0(N5723));
MXI2XL addgen2_A_I1262 (.Y(N692), .A(N5732), .B(N5729), .S0(N3097));
MXI2X1 addgen2_A_I1263 (.Y(N3106), .A(N5631), .B(N5630), .S0(N5723));
MXI2X1 addgen2_A_I1264 (.Y(N693), .A(N5732), .B(N5729), .S0(N3106));
MXI2XL addgen2_A_I1265 (.Y(N3115), .A(N5632), .B(N5631), .S0(N5723));
MXI2XL addgen2_A_I1266 (.Y(N694), .A(N5732), .B(N5729), .S0(N3115));
MXI2XL addgen2_A_I1267 (.Y(N3124), .A(N5633), .B(N5632), .S0(N5723));
MXI2XL addgen2_A_I1268 (.Y(N695), .A(N5732), .B(N5729), .S0(N3124));
MXI2XL addgen2_A_I1269 (.Y(N3133), .A(N5634), .B(N5633), .S0(N5723));
MXI2XL addgen2_A_I1270 (.Y(N696), .A(N5732), .B(N5729), .S0(N3133));
MXI2XL addgen2_A_I1271 (.Y(N3142), .A(N5635), .B(N5634), .S0(N5723));
MXI2XL addgen2_A_I1272 (.Y(N697), .A(N5732), .B(N5729), .S0(N3142));
MXI2XL addgen2_A_I1273 (.Y(N3151), .A(N5636), .B(N5635), .S0(N5723));
MXI2XL addgen2_A_I1274 (.Y(N698), .A(N5732), .B(N5731), .S0(N3151));
MXI2XL addgen2_A_I1275 (.Y(N3160), .A(N5637), .B(N5636), .S0(N5723));
MXI2XL addgen2_A_I1276 (.Y(N699), .A(N5732), .B(N5731), .S0(N3160));
MXI2XL addgen2_A_I1277 (.Y(N3169), .A(N5638), .B(N5637), .S0(N5723));
MXI2XL addgen2_A_I1278 (.Y(N700), .A(N5732), .B(N5731), .S0(N3169));
MXI2XL addgen2_A_I1279 (.Y(N3178), .A(N5639), .B(N5638), .S0(N5723));
MXI2XL addgen2_A_I1280 (.Y(N701), .A(N5732), .B(N5731), .S0(N3178));
MXI2XL addgen2_A_I1281 (.Y(N3187), .A(N5640), .B(N5639), .S0(N5723));
MXI2XL addgen2_A_I1282 (.Y(N702), .A(N5732), .B(N5731), .S0(N3187));
MXI2XL addgen2_A_I1283 (.Y(N3196), .A(N5641), .B(N5640), .S0(N5723));
MXI2XL addgen2_A_I1284 (.Y(N703), .A(N5732), .B(N5731), .S0(N3196));
MXI2XL addgen2_A_I1285 (.Y(N3205), .A(N5642), .B(N5641), .S0(N5723));
MXI2XL addgen2_A_I1286 (.Y(N704), .A(N5732), .B(N5731), .S0(N3205));
NAND2XL addgen2_A_I1287 (.Y(N3214), .A(N5642), .B(N5723));
MXI2XL addgen2_A_I1288 (.Y(N705), .A(N5732), .B(N5731), .S0(N3214));
XNOR2X1 enc2_A_I1289 (.Y(N709), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
NAND2XL enc2_A_I1290 (.Y(N3223), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
NOR2XL enc2_A_I1291 (.Y(N3225), .A(inst_cellmath__203_0_in1[28]), .B(inst_cellmath__203_0_in1[27]));
AND2XL enc2_A_I1292 (.Y(N711), .A(N3223), .B(inst_cellmath__203_0_in1[29]));
NOR2XL enc2_A_I1293 (.Y(N710), .A(N3225), .B(inst_cellmath__203_0_in1[29]));
INVX2 inst_cellmath__203_0_I1935 (.Y(N5733), .A(N709));
INVXL inst_cellmath__203_0_I1941 (.Y(N5739), .A(N5733));
INVX2 inst_cellmath__203_0_I1940 (.Y(N5738), .A(N5733));
INVX2 inst_cellmath__203_0_I1939 (.Y(N5737), .A(N5733));
INVXL inst_cellmath__203_0_I1938 (.Y(N5736), .A(N5733));
INVXL inst_cellmath__203_0_I1949 (.Y(N5747), .A(N710));
INVXL inst_cellmath__203_0_I1947 (.Y(N5745), .A(N710));
INVX1 inst_cellmath__203_0_I1950 (.Y(N5748), .A(N711));
NOR2XL addgen2_A_I1294 (.Y(N3236), .A(N5617), .B(N5738));
MXI2XL addgen2_A_I1295 (.Y(N715), .A(N5748), .B(N5747), .S0(N3236));
MXI2XL addgen2_A_I1296 (.Y(N3245), .A(N5624), .B(N5617), .S0(N5739));
MXI2XL addgen2_A_I1297 (.Y(N716), .A(N5748), .B(N5747), .S0(N3245));
MXI2XL addgen2_A_I1298 (.Y(N3254), .A(N5625), .B(N5624), .S0(N5738));
MXI2XL addgen2_A_I1299 (.Y(N717), .A(N5748), .B(N5747), .S0(N3254));
MXI2XL addgen2_A_I1300 (.Y(N3263), .A(N5626), .B(N5625), .S0(N5738));
MXI2XL addgen2_A_I1301 (.Y(N718), .A(N5748), .B(N5747), .S0(N3263));
MXI2XL addgen2_A_I1302 (.Y(N3272), .A(N5627), .B(N5626), .S0(N5738));
MXI2XL addgen2_A_I1303 (.Y(N719), .A(N5748), .B(N5747), .S0(N3272));
MXI2XL addgen2_A_I1304 (.Y(N3281), .A(N5628), .B(N5627), .S0(N5738));
MXI2XL addgen2_A_I1305 (.Y(N720), .A(N5748), .B(N5745), .S0(N3281));
MXI2XL addgen2_A_I1306 (.Y(N3290), .A(N5629), .B(N5628), .S0(N5737));
MXI2XL addgen2_A_I1307 (.Y(N721), .A(N5748), .B(N5745), .S0(N3290));
MXI2XL addgen2_A_I1308 (.Y(N3299), .A(N5630), .B(N5629), .S0(N5737));
MXI2XL addgen2_A_I1309 (.Y(N722), .A(N5748), .B(N5745), .S0(N3299));
MXI2XL addgen2_A_I1310 (.Y(N3308), .A(N5631), .B(N5630), .S0(N5737));
MXI2XL addgen2_A_I1311 (.Y(N723), .A(N5748), .B(N5745), .S0(N3308));
MXI2XL addgen2_A_I1312 (.Y(N3317), .A(N5632), .B(N5631), .S0(N5737));
MXI2XL addgen2_A_I1313 (.Y(N724), .A(N5748), .B(N5745), .S0(N3317));
MXI2XL addgen2_A_I1314 (.Y(N3326), .A(N5633), .B(N5632), .S0(N5736));
MXI2XL addgen2_A_I1315 (.Y(N725), .A(N5748), .B(N5745), .S0(N3326));
MXI2XL addgen2_A_I1316 (.Y(N3335), .A(N5634), .B(N5633), .S0(N5736));
MXI2XL addgen2_A_I1317 (.Y(N726), .A(N5748), .B(N5745), .S0(N3335));
MXI2XL addgen2_A_I1318 (.Y(N3344), .A(N5635), .B(N5634), .S0(N5736));
MXI2XL addgen2_A_I1319 (.Y(N727), .A(N5748), .B(N5745), .S0(N3344));
MXI2XL addgen2_A_I1320 (.Y(N3353), .A(N5636), .B(N5635), .S0(N5736));
MXI2XL addgen2_A_I1321 (.Y(N728), .A(N5748), .B(N5747), .S0(N3353));
MXI2XL addgen2_A_I1322 (.Y(N3362), .A(N5637), .B(N5636), .S0(N5739));
MXI2XL addgen2_A_I1323 (.Y(N729), .A(N5748), .B(N5747), .S0(N3362));
MXI2XL addgen2_A_I1324 (.Y(N3371), .A(N5638), .B(N5637), .S0(N5739));
MXI2XL addgen2_A_I1325 (.Y(N730), .A(N5748), .B(N5747), .S0(N3371));
MXI2XL addgen2_A_I1326 (.Y(N3380), .A(N5639), .B(N5638), .S0(N5739));
MXI2XL addgen2_A_I1327 (.Y(N731), .A(N5748), .B(N5747), .S0(N3380));
MXI2XL addgen2_A_I1328 (.Y(N3389), .A(N5640), .B(N5639), .S0(N5739));
MXI2XL addgen2_A_I1329 (.Y(N732), .A(N5748), .B(N5747), .S0(N3389));
MXI2XL addgen2_A_I1330 (.Y(N3398), .A(N5641), .B(N5640), .S0(N5738));
MXI2XL addgen2_A_I1331 (.Y(N733), .A(N5748), .B(N5747), .S0(N3398));
MXI2XL addgen2_A_I1332 (.Y(N3407), .A(N5642), .B(N5641), .S0(N5738));
MXI2XL addgen2_A_I1333 (.Y(N734), .A(N5748), .B(N5747), .S0(N3407));
NAND2XL addgen2_A_I1334 (.Y(N3416), .A(N5642), .B(N5738));
MXI2XL addgen2_A_I1335 (.Y(N735), .A(N5748), .B(N5747), .S0(N3416));
NAND2XL enc2_A_I1337 (.Y(N3425), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
NOR2XL enc2_A_I1338 (.Y(N3427), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
AND2XL enc2_A_I1339 (.Y(N741), .A(N3425), .B(inst_cellmath__203_0_in1[31]));
XOR2XL inst_cellmath__203_0_I2218 (.Y(N5749), .A(inst_cellmath__203_0_in1[30]), .B(inst_cellmath__203_0_in1[29]));
INVXL inst_cellmath__203_0_I1957 (.Y(N5755), .A(N5749));
INVX2 inst_cellmath__203_0_I1956 (.Y(N5754), .A(N5749));
OR2X1 inst_cellmath__203_0_I2219 (.Y(N5763), .A(N3427), .B(inst_cellmath__203_0_in1[31]));
INVX1 inst_cellmath__203_0_I1966 (.Y(N5764), .A(N741));
NOR2XL addgen2_A_I1341 (.Y(N3438), .A(N5617), .B(N5754));
MXI2XL addgen2_A_I1342 (.Y(N745), .A(N5764), .B(N5763), .S0(N3438));
MXI2XL addgen2_A_I1343 (.Y(N3447), .A(N5624), .B(N5617), .S0(N5755));
MXI2XL addgen2_A_I1344 (.Y(N746), .A(N5764), .B(N5763), .S0(N3447));
MXI2XL addgen2_A_I1345 (.Y(N3456), .A(N5625), .B(N5624), .S0(N5754));
MXI2XL addgen2_A_I1346 (.Y(N747), .A(N5764), .B(N5763), .S0(N3456));
MXI2XL addgen2_A_I1347 (.Y(N3465), .A(N5626), .B(N5625), .S0(N5754));
MXI2XL addgen2_A_I1348 (.Y(N748), .A(N5764), .B(N5763), .S0(N3465));
MXI2XL addgen2_A_I1349 (.Y(N3474), .A(N5627), .B(N5626), .S0(N5754));
MXI2XL addgen2_A_I1350 (.Y(N749), .A(N5764), .B(N5763), .S0(N3474));
MXI2XL addgen2_A_I1351 (.Y(N3483), .A(N5628), .B(N5627), .S0(N5754));
MXI2XL addgen2_A_I1352 (.Y(N750), .A(N5764), .B(N5763), .S0(N3483));
MXI2XL addgen2_A_I1353 (.Y(N3492), .A(N5629), .B(N5628), .S0(N5754));
MXI2XL addgen2_A_I1354 (.Y(N751), .A(N5764), .B(N5763), .S0(N3492));
MXI2XL addgen2_A_I1355 (.Y(N3501), .A(N5630), .B(N5629), .S0(N5754));
MXI2XL addgen2_A_I1356 (.Y(N752), .A(N5764), .B(N5763), .S0(N3501));
MXI2XL addgen2_A_I1357 (.Y(N3510), .A(N5631), .B(N5630), .S0(N5754));
MXI2XL addgen2_A_I1358 (.Y(N753), .A(N5764), .B(N5763), .S0(N3510));
MXI2XL addgen2_A_I1359 (.Y(N3519), .A(N5632), .B(N5631), .S0(N5754));
MXI2XL addgen2_A_I1360 (.Y(N754), .A(N5764), .B(N5763), .S0(N3519));
MXI2XL addgen2_A_I1361 (.Y(N3528), .A(N5633), .B(N5632), .S0(N5754));
MXI2XL addgen2_A_I1362 (.Y(N755), .A(N5764), .B(N5763), .S0(N3528));
MXI2XL addgen2_A_I1363 (.Y(N3537), .A(N5634), .B(N5633), .S0(N5754));
MXI2XL addgen2_A_I1364 (.Y(N756), .A(N5764), .B(N5763), .S0(N3537));
MXI2XL addgen2_A_I1365 (.Y(N3546), .A(N5635), .B(N5634), .S0(N5754));
MXI2XL addgen2_A_I1366 (.Y(N757), .A(N5764), .B(N5763), .S0(N3546));
MXI2XL addgen2_A_I1367 (.Y(N3555), .A(N5636), .B(N5635), .S0(N5754));
MXI2XL addgen2_A_I1368 (.Y(N758), .A(N5764), .B(N5763), .S0(N3555));
MXI2XL addgen2_A_I1369 (.Y(N3564), .A(N5637), .B(N5636), .S0(N5755));
MXI2XL addgen2_A_I1370 (.Y(N759), .A(N5764), .B(N5763), .S0(N3564));
MXI2XL addgen2_A_I1371 (.Y(N3573), .A(N5638), .B(N5637), .S0(N5755));
MXI2XL addgen2_A_I1372 (.Y(N760), .A(N5764), .B(N5763), .S0(N3573));
MXI2XL addgen2_A_I1373 (.Y(N3582), .A(N5639), .B(N5638), .S0(N5755));
MXI2XL addgen2_A_I1374 (.Y(N761), .A(N5764), .B(N5763), .S0(N3582));
MXI2XL addgen2_A_I1375 (.Y(N3591), .A(N5640), .B(N5639), .S0(N5755));
MXI2XL addgen2_A_I1376 (.Y(N762), .A(N5764), .B(N5763), .S0(N3591));
MXI2XL addgen2_A_I1377 (.Y(N3600), .A(N5641), .B(N5640), .S0(N5754));
MXI2XL addgen2_A_I1378 (.Y(N763), .A(N5764), .B(N5763), .S0(N3600));
MXI2XL addgen2_A_I1379 (.Y(N3609), .A(N5642), .B(N5641), .S0(N5754));
MXI2XL addgen2_A_I1380 (.Y(N764), .A(N5764), .B(N5763), .S0(N3609));
NAND2XL addgen2_A_I1381 (.Y(N3618), .A(N5642), .B(N5754));
MXI2XL addgen2_A_I1382 (.Y(N765), .A(N5764), .B(N5763), .S0(N3618));
ADDHX1 inst_cellmath__203_0_I281 (.CO(N770), .S(N768), .A(inst_cellmath__203_0_in1[32]), .B(inst_cellmath__203_0_in1[31]));
INVX3 inst_cellmath__203_0_I1967 (.Y(N5765), .A(N768));
INVX2 inst_cellmath__203_0_I1968 (.Y(N5766), .A(N770));
NOR2XL inst_cellmath__203_0_I285 (.Y(N779), .A(N5765), .B(N5617));
OAI22XL inst_cellmath__203_0_I286 (.Y(N781), .A0(N5617), .A1(N5766), .B0(N5765), .B1(N5624));
OAI22XL inst_cellmath__203_0_I287 (.Y(N783), .A0(N5624), .A1(N5766), .B0(N5765), .B1(N5625));
OAI22XL inst_cellmath__203_0_I288 (.Y(N785), .A0(N5625), .A1(N5766), .B0(N5765), .B1(N5626));
OAI22XL inst_cellmath__203_0_I289 (.Y(N787), .A0(N5626), .A1(N5766), .B0(N5765), .B1(N5627));
OAI22XL inst_cellmath__203_0_I290 (.Y(N789), .A0(N5627), .A1(N5766), .B0(N5765), .B1(N5628));
OAI22XL inst_cellmath__203_0_I291 (.Y(N791), .A0(N5628), .A1(N5766), .B0(N5765), .B1(N5629));
OAI22XL inst_cellmath__203_0_I292 (.Y(N793), .A0(N5629), .A1(N5766), .B0(N5765), .B1(N5630));
OAI22XL inst_cellmath__203_0_I293 (.Y(N795), .A0(N5630), .A1(N5766), .B0(N5765), .B1(N5631));
OAI22XL inst_cellmath__203_0_I294 (.Y(N797), .A0(N5631), .A1(N5766), .B0(N5765), .B1(N5632));
OAI22XL inst_cellmath__203_0_I295 (.Y(N799), .A0(N5632), .A1(N5766), .B0(N5765), .B1(N5633));
OAI22XL inst_cellmath__203_0_I296 (.Y(N801), .A0(N5633), .A1(N5766), .B0(N5765), .B1(N5634));
OAI22XL inst_cellmath__203_0_I297 (.Y(N803), .A0(N5634), .A1(N5766), .B0(N5765), .B1(N5635));
OAI22XL inst_cellmath__203_0_I298 (.Y(N805), .A0(N5635), .A1(N5766), .B0(N5765), .B1(N5636));
OAI22XL inst_cellmath__203_0_I299 (.Y(N807), .A0(N5636), .A1(N5766), .B0(N5765), .B1(N5637));
OAI22XL inst_cellmath__203_0_I300 (.Y(N809), .A0(N5637), .A1(N5766), .B0(N5765), .B1(N5638));
OAI22XL inst_cellmath__203_0_I301 (.Y(N811), .A0(N5638), .A1(N5766), .B0(N5765), .B1(N5639));
OAI22XL inst_cellmath__203_0_I302 (.Y(N813), .A0(N5639), .A1(N5766), .B0(N5765), .B1(N5640));
OAI22XL inst_cellmath__203_0_I303 (.Y(N815), .A0(N5640), .A1(N5766), .B0(N5765), .B1(N5641));
OAI22XL inst_cellmath__203_0_I304 (.Y(N817), .A0(N5641), .A1(N5766), .B0(N5765), .B1(N5642));
OAI21XL inst_cellmath__203_0_I305 (.Y(N819), .A0(N5766), .A1(N5642), .B0(N5765));
AND2XL inst_cellmath__203_0_I306 (.Y(N1366), .A(N5766), .B(N5765));
INVX1 inst_cellmath__203_0_I1969 (.Y(N5767), .A(inst_cellmath__203_0_in3[0]));
INVX2 inst_cellmath__203_0_I1970 (.Y(N5768), .A(inst_cellmath__203_0_in3[1]));
INVX1 inst_cellmath__203_0_I1971 (.Y(N5769), .A(inst_cellmath__203_0_in3[2]));
INVX2 inst_cellmath__203_0_I1972 (.Y(N5770), .A(inst_cellmath__203_0_in3[3]));
INVX2 inst_cellmath__203_0_I1973 (.Y(N5771), .A(inst_cellmath__203_0_in3[4]));
INVX2 inst_cellmath__203_0_I1974 (.Y(N5772), .A(inst_cellmath__203_0_in3[5]));
INVX2 inst_cellmath__203_0_I1975 (.Y(N5773), .A(inst_cellmath__203_0_in3[6]));
INVX2 inst_cellmath__203_0_I1976 (.Y(N5774), .A(inst_cellmath__203_0_in3[7]));
INVX2 inst_cellmath__203_0_I1977 (.Y(N5775), .A(inst_cellmath__203_0_in3[8]));
INVX1 inst_cellmath__203_0_I1978 (.Y(N5776), .A(inst_cellmath__203_0_in3[9]));
INVX2 inst_cellmath__203_0_I1979 (.Y(N5777), .A(inst_cellmath__203_0_in3[10]));
INVX1 inst_cellmath__203_0_I1980 (.Y(N5778), .A(inst_cellmath__203_0_in3[11]));
INVX2 inst_cellmath__203_0_I1981 (.Y(N5779), .A(inst_cellmath__203_0_in3[12]));
INVX2 inst_cellmath__203_0_I1982 (.Y(N5780), .A(inst_cellmath__203_0_in3[13]));
INVX1 inst_cellmath__203_0_I1983 (.Y(N5781), .A(inst_cellmath__203_0_in3[14]));
INVX1 inst_cellmath__203_0_I1984 (.Y(N5782), .A(inst_cellmath__203_0_in3[15]));
INVX2 inst_cellmath__203_0_I1985 (.Y(N5783), .A(inst_cellmath__203_0_in3[16]));
INVX1 inst_cellmath__203_0_I1986 (.Y(N5784), .A(inst_cellmath__203_0_in3[17]));
INVX1 inst_cellmath__203_0_I1987 (.Y(N5785), .A(inst_cellmath__203_0_in3[18]));
INVXL inst_cellmath__203_0_I1988 (.Y(N5786), .A(inst_cellmath__203_0_in3[19]));
INVXL inst_cellmath__203_0_I1989 (.Y(N5787), .A(inst_cellmath__203_0_in3[20]));
INVXL inst_cellmath__203_0_I1990 (.Y(N5788), .A(inst_cellmath__203_0_in3[21]));
INVXL inst_cellmath__203_0_I1991 (.Y(N5789), .A(inst_cellmath__203_0_in0[0]));
NOR2XL inst_cellmath__203_0_I382 (.Y(N1025), .A(N5789), .B(N5767));
NOR2XL inst_cellmath__203_0_I383 (.Y(N1027), .A(N5789), .B(N5768));
NOR2XL inst_cellmath__203_0_I384 (.Y(N1029), .A(N5789), .B(N5769));
NOR2XL inst_cellmath__203_0_I385 (.Y(N1031), .A(N5789), .B(N5770));
NOR2XL inst_cellmath__203_0_I386 (.Y(N1033), .A(N5789), .B(N5771));
NOR2XL inst_cellmath__203_0_I387 (.Y(N1035), .A(N5789), .B(N5772));
NOR2XL inst_cellmath__203_0_I388 (.Y(N1037), .A(N5789), .B(N5773));
NOR2XL inst_cellmath__203_0_I389 (.Y(N1039), .A(N5789), .B(N5774));
NOR2XL inst_cellmath__203_0_I390 (.Y(N1041), .A(N5789), .B(N5775));
NOR2XL inst_cellmath__203_0_I391 (.Y(N1043), .A(N5789), .B(N5776));
NOR2XL inst_cellmath__203_0_I392 (.Y(N1045), .A(N5789), .B(N5777));
NOR2XL inst_cellmath__203_0_I393 (.Y(N1047), .A(N5789), .B(N5778));
NOR2XL inst_cellmath__203_0_I394 (.Y(N1049), .A(N5789), .B(N5779));
NOR2XL inst_cellmath__203_0_I395 (.Y(N1051), .A(N5789), .B(N5780));
NOR2XL inst_cellmath__203_0_I396 (.Y(N1053), .A(N5789), .B(N5781));
NOR2XL inst_cellmath__203_0_I397 (.Y(N1055), .A(N5789), .B(N5782));
NOR2XL inst_cellmath__203_0_I398 (.Y(N1698), .A(N5789), .B(N5783));
NOR2XL inst_cellmath__203_0_I399 (.Y(N1732), .A(N5789), .B(N5784));
NOR2XL inst_cellmath__203_0_I400 (.Y(N1061), .A(N5789), .B(N5785));
NOR2XL inst_cellmath__203_0_I401 (.Y(N1798), .A(N5789), .B(N5786));
NOR2XL inst_cellmath__203_0_I402 (.Y(N1830), .A(N5789), .B(N5787));
NOR2XL inst_cellmath__203_0_I403 (.Y(N1067), .A(N5789), .B(N5788));
INVXL inst_cellmath__203_0_I1999 (.Y(N5797), .A(inst_cellmath__203_0_in0[1]));
NAND2BX1 inst_cellmath__203_0_I2220 (.Y(N5805), .AN(inst_cellmath__203_0_in0[2]), .B(inst_cellmath__203_0_in0[1]));
INVXL inst_cellmath__203_0_I2008 (.Y(N5806), .A(inst_cellmath__203_0_in0[2]));
NOR2XL addgen2_A_I1388 (.Y(N3640), .A(N5767), .B(N5797));
MXI2XL addgen2_A_I1389 (.Y(N1077), .A(N5806), .B(N5805), .S0(N3640));
MXI2XL addgen2_A_I1390 (.Y(N3649), .A(N5768), .B(N5767), .S0(N5797));
MXI2XL addgen2_A_I1391 (.Y(N1078), .A(N5806), .B(N5805), .S0(N3649));
MXI2XL addgen2_A_I1392 (.Y(N3658), .A(N5769), .B(N5768), .S0(N5797));
MXI2XL addgen2_A_I1393 (.Y(N1079), .A(N5806), .B(N5805), .S0(N3658));
MXI2XL addgen2_A_I1394 (.Y(N3667), .A(N5770), .B(N5769), .S0(N5797));
MXI2XL addgen2_A_I1395 (.Y(N1080), .A(N5806), .B(N5805), .S0(N3667));
MXI2XL addgen2_A_I1396 (.Y(N3676), .A(N5771), .B(N5770), .S0(N5797));
MXI2XL addgen2_A_I1397 (.Y(N1081), .A(N5806), .B(N5805), .S0(N3676));
MXI2XL addgen2_A_I1398 (.Y(N3685), .A(N5772), .B(N5771), .S0(N5797));
MXI2XL addgen2_A_I1399 (.Y(N1082), .A(N5806), .B(N5805), .S0(N3685));
MXI2XL addgen2_A_I1400 (.Y(N3694), .A(N5773), .B(N5772), .S0(N5797));
MXI2XL addgen2_A_I1401 (.Y(N1083), .A(N5806), .B(N5805), .S0(N3694));
MXI2XL addgen2_A_I1402 (.Y(N3703), .A(N5774), .B(N5773), .S0(N5797));
MXI2XL addgen2_A_I1403 (.Y(N1084), .A(N5806), .B(N5805), .S0(N3703));
MXI2XL addgen2_A_I1404 (.Y(N3712), .A(N5775), .B(N5774), .S0(N5797));
MXI2XL addgen2_A_I1405 (.Y(N1085), .A(N5806), .B(N5805), .S0(N3712));
MXI2XL addgen2_A_I1406 (.Y(N3721), .A(N5776), .B(N5775), .S0(N5797));
MXI2XL addgen2_A_I1407 (.Y(N1086), .A(N5806), .B(N5805), .S0(N3721));
MXI2XL addgen2_A_I1408 (.Y(N3730), .A(N5777), .B(N5776), .S0(N5797));
MXI2XL addgen2_A_I1409 (.Y(N1087), .A(N5806), .B(N5805), .S0(N3730));
MXI2XL addgen2_A_I1410 (.Y(N3739), .A(N5778), .B(N5777), .S0(N5797));
MXI2XL addgen2_A_I1411 (.Y(N1088), .A(N5806), .B(N5805), .S0(N3739));
MXI2XL addgen2_A_I1412 (.Y(N3748), .A(N5779), .B(N5778), .S0(N5797));
MXI2XL addgen2_A_I1413 (.Y(N1089), .A(N5806), .B(N5805), .S0(N3748));
MXI2XL addgen2_A_I1414 (.Y(N3757), .A(N5780), .B(N5779), .S0(N5797));
MXI2XL addgen2_A_I1415 (.Y(N1090), .A(N5806), .B(N5805), .S0(N3757));
MXI2XL addgen2_A_I1416 (.Y(N3766), .A(N5781), .B(N5780), .S0(N5797));
MXI2XL addgen2_A_I1417 (.Y(N1091), .A(N5806), .B(N5805), .S0(N3766));
MXI2XL addgen2_A_I1418 (.Y(N3775), .A(N5782), .B(N5781), .S0(N5797));
MXI2XL addgen2_A_I1419 (.Y(N1092), .A(N5806), .B(N5805), .S0(N3775));
MXI2XL addgen2_A_I1420 (.Y(N3784), .A(N5783), .B(N5782), .S0(N5797));
MXI2XL addgen2_A_I1421 (.Y(N1093), .A(N5806), .B(N5805), .S0(N3784));
MXI2XL addgen2_A_I1422 (.Y(N3793), .A(N5784), .B(N5783), .S0(N5797));
MXI2XL addgen2_A_I1423 (.Y(N1094), .A(N5806), .B(N5805), .S0(N3793));
MXI2XL addgen2_A_I1424 (.Y(N3802), .A(N5785), .B(N5784), .S0(N5797));
MXI2XL addgen2_A_I1425 (.Y(N1095), .A(N5806), .B(N5805), .S0(N3802));
MXI2XL addgen2_A_I1426 (.Y(N3811), .A(N5786), .B(N5785), .S0(N5797));
MXI2XL addgen2_A_I1427 (.Y(N1096), .A(N5806), .B(N5805), .S0(N3811));
MXI2XL addgen2_A_I1428 (.Y(N3820), .A(N5787), .B(N5786), .S0(N5797));
MXI2XL addgen2_A_I1429 (.Y(N1097), .A(N5806), .B(N5805), .S0(N3820));
MXI2XL addgen2_A_I1430 (.Y(N3829), .A(N5788), .B(N5787), .S0(N5797));
MXI2XL addgen2_A_I1431 (.Y(N1098), .A(N5806), .B(N5805), .S0(N3829));
NOR2BX1 addgen2_A_I1432 (.Y(N3838), .AN(N5797), .B(N5788));
MXI2XL addgen2_A_I1433 (.Y(N1099), .A(N5806), .B(N5805), .S0(N3838));
CLKINVX1 inst_cellmath__203_0_I2017 (.Y(N5815), .A(inst_cellmath__203_0_in0[3]));
INVXL inst_cellmath__203_0_I2018 (.Y(N5816), .A(N5815));
XNOR2X1 enc2_A_I1434 (.Y(N1103), .A(N5816), .B(inst_cellmath__203_0_in0[2]));
NAND2XL enc2_A_I1435 (.Y(N3847), .A(N5816), .B(inst_cellmath__203_0_in0[2]));
NOR2XL enc2_A_I1436 (.Y(N3849), .A(N5816), .B(inst_cellmath__203_0_in0[2]));
CLKINVX1 inst_cellmath__203_0_I2019 (.Y(N5817), .A(inst_cellmath__203_0_in0[4]));
INVXL inst_cellmath__203_0_I2020 (.Y(N5818), .A(N5817));
AND2XL enc2_A_I1437 (.Y(N1105), .A(N3847), .B(N5818));
OR2XL inst_cellmath__203_0_I2223 (.Y(N5833), .A(N3849), .B(N5818));
INVXL inst_cellmath__203_0_I2044 (.Y(N5842), .A(N1105));
NOR2XL addgen2_A_I1439 (.Y(N3860), .A(N5767), .B(N1103));
MXI2XL addgen2_A_I1440 (.Y(N1109), .A(N5842), .B(N5833), .S0(N3860));
MXI2XL addgen2_A_I1441 (.Y(N3869), .A(N5768), .B(N5767), .S0(N1103));
MXI2XL addgen2_A_I1442 (.Y(N1110), .A(N5842), .B(N5833), .S0(N3869));
MXI2XL addgen2_A_I1443 (.Y(N3878), .A(N5769), .B(N5768), .S0(N1103));
MXI2XL addgen2_A_I1444 (.Y(N1111), .A(N5842), .B(N5833), .S0(N3878));
MXI2XL addgen2_A_I1445 (.Y(N3887), .A(N5770), .B(N5769), .S0(N1103));
MXI2XL addgen2_A_I1446 (.Y(N1112), .A(N5842), .B(N5833), .S0(N3887));
MXI2XL addgen2_A_I1447 (.Y(N3896), .A(N5771), .B(N5770), .S0(N1103));
MXI2XL addgen2_A_I1448 (.Y(N1113), .A(N5842), .B(N5833), .S0(N3896));
MXI2XL addgen2_A_I1449 (.Y(N3905), .A(N5772), .B(N5771), .S0(N1103));
MXI2XL addgen2_A_I1450 (.Y(N1114), .A(N5842), .B(N5833), .S0(N3905));
MXI2XL addgen2_A_I1451 (.Y(N3914), .A(N5773), .B(N5772), .S0(N1103));
MXI2XL addgen2_A_I1452 (.Y(N1115), .A(N5842), .B(N5833), .S0(N3914));
MXI2XL addgen2_A_I1453 (.Y(N3923), .A(N5774), .B(N5773), .S0(N1103));
MXI2XL addgen2_A_I1454 (.Y(N1116), .A(N5842), .B(N5833), .S0(N3923));
MXI2XL addgen2_A_I1455 (.Y(N3932), .A(N5775), .B(N5774), .S0(N1103));
MXI2XL addgen2_A_I1456 (.Y(N1117), .A(N5842), .B(N5833), .S0(N3932));
MXI2XL addgen2_A_I1457 (.Y(N3941), .A(N5776), .B(N5775), .S0(N1103));
MXI2XL addgen2_A_I1458 (.Y(N1118), .A(N5842), .B(N5833), .S0(N3941));
MXI2XL addgen2_A_I1459 (.Y(N3950), .A(N5777), .B(N5776), .S0(N1103));
MXI2XL addgen2_A_I1460 (.Y(N1119), .A(N5842), .B(N5833), .S0(N3950));
MXI2XL addgen2_A_I1461 (.Y(N3959), .A(N5778), .B(N5777), .S0(N1103));
MXI2XL addgen2_A_I1462 (.Y(N1120), .A(N5842), .B(N5833), .S0(N3959));
MXI2XL addgen2_A_I1463 (.Y(N3968), .A(N5779), .B(N5778), .S0(N1103));
MXI2XL addgen2_A_I1464 (.Y(N1121), .A(N5842), .B(N5833), .S0(N3968));
MXI2XL addgen2_A_I1465 (.Y(N3977), .A(N5780), .B(N5779), .S0(N1103));
MXI2XL addgen2_A_I1466 (.Y(N1122), .A(N5842), .B(N5833), .S0(N3977));
MXI2XL addgen2_A_I1467 (.Y(N3986), .A(N5781), .B(N5780), .S0(N1103));
MXI2XL addgen2_A_I1468 (.Y(N1123), .A(N5842), .B(N5833), .S0(N3986));
MXI2XL addgen2_A_I1469 (.Y(N3995), .A(N5782), .B(N5781), .S0(N1103));
MXI2XL addgen2_A_I1470 (.Y(N1124), .A(N5842), .B(N5833), .S0(N3995));
MXI2XL addgen2_A_I1471 (.Y(N4004), .A(N5783), .B(N5782), .S0(N1103));
MXI2XL addgen2_A_I1472 (.Y(N1125), .A(N5842), .B(N5833), .S0(N4004));
MXI2XL addgen2_A_I1473 (.Y(N4013), .A(N5784), .B(N5783), .S0(N1103));
MXI2XL addgen2_A_I1474 (.Y(N1126), .A(N5842), .B(N5833), .S0(N4013));
MXI2XL addgen2_A_I1475 (.Y(N4022), .A(N5785), .B(N5784), .S0(N1103));
MXI2XL addgen2_A_I1476 (.Y(N1127), .A(N5842), .B(N5833), .S0(N4022));
MXI2XL addgen2_A_I1477 (.Y(N4031), .A(N5786), .B(N5785), .S0(N1103));
MXI2XL addgen2_A_I1478 (.Y(N1128), .A(N5842), .B(N5833), .S0(N4031));
MXI2XL addgen2_A_I1479 (.Y(N4040), .A(N5787), .B(N5786), .S0(N1103));
MXI2XL addgen2_A_I1480 (.Y(N1129), .A(N5842), .B(N5833), .S0(N4040));
MXI2XL addgen2_A_I1481 (.Y(N4049), .A(N5788), .B(N5787), .S0(N1103));
MXI2XL addgen2_A_I1482 (.Y(N1130), .A(N5842), .B(N5833), .S0(N4049));
NOR2BX1 addgen2_A_I1483 (.Y(N4058), .AN(N1103), .B(N5788));
MXI2XL addgen2_A_I1484 (.Y(N1131), .A(N5842), .B(N5833), .S0(N4058));
XNOR2X1 enc2_A_I1485 (.Y(N1135), .A(inst_cellmath__203_0_in0[5]), .B(N5818));
NAND2XL enc2_A_I1486 (.Y(N4067), .A(inst_cellmath__203_0_in0[5]), .B(N5818));
NOR2XL enc2_A_I1487 (.Y(N4069), .A(inst_cellmath__203_0_in0[5]), .B(N5818));
CLKINVX1 inst_cellmath__203_0_I2045 (.Y(N5843), .A(inst_cellmath__203_0_in0[6]));
INVXL inst_cellmath__203_0_I2046 (.Y(N5844), .A(N5843));
AND2XL enc2_A_I1488 (.Y(N1137), .A(N4067), .B(N5844));
OR2XL inst_cellmath__203_0_I2225 (.Y(N5859), .A(N4069), .B(N5844));
INVXL inst_cellmath__203_0_I2070 (.Y(N5868), .A(N1137));
NOR2XL addgen2_A_I1490 (.Y(N4080), .A(N5767), .B(N1135));
MXI2XL addgen2_A_I1491 (.Y(N1141), .A(N5868), .B(N5859), .S0(N4080));
MXI2XL addgen2_A_I1492 (.Y(N4089), .A(N5768), .B(N5767), .S0(N1135));
MXI2XL addgen2_A_I1493 (.Y(N1142), .A(N5868), .B(N5859), .S0(N4089));
MXI2XL addgen2_A_I1494 (.Y(N4098), .A(N5769), .B(N5768), .S0(N1135));
MXI2XL addgen2_A_I1495 (.Y(N1143), .A(N5868), .B(N5859), .S0(N4098));
MXI2XL addgen2_A_I1496 (.Y(N4107), .A(N5770), .B(N5769), .S0(N1135));
MXI2XL addgen2_A_I1497 (.Y(N1144), .A(N5868), .B(N5859), .S0(N4107));
MXI2XL addgen2_A_I1498 (.Y(N4116), .A(N5771), .B(N5770), .S0(N1135));
MXI2XL addgen2_A_I1499 (.Y(N1145), .A(N5868), .B(N5859), .S0(N4116));
MXI2XL addgen2_A_I1500 (.Y(N4125), .A(N5772), .B(N5771), .S0(N1135));
MXI2XL addgen2_A_I1501 (.Y(N1146), .A(N5868), .B(N5859), .S0(N4125));
MXI2XL addgen2_A_I1502 (.Y(N4134), .A(N5773), .B(N5772), .S0(N1135));
MXI2XL addgen2_A_I1503 (.Y(N1147), .A(N5868), .B(N5859), .S0(N4134));
MXI2XL addgen2_A_I1504 (.Y(N4143), .A(N5774), .B(N5773), .S0(N1135));
MXI2XL addgen2_A_I1505 (.Y(N1148), .A(N5868), .B(N5859), .S0(N4143));
MXI2XL addgen2_A_I1506 (.Y(N4152), .A(N5775), .B(N5774), .S0(N1135));
MXI2XL addgen2_A_I1507 (.Y(N1149), .A(N5868), .B(N5859), .S0(N4152));
MXI2XL addgen2_A_I1508 (.Y(N4161), .A(N5776), .B(N5775), .S0(N1135));
MXI2XL addgen2_A_I1509 (.Y(N1150), .A(N5868), .B(N5859), .S0(N4161));
MXI2XL addgen2_A_I1510 (.Y(N4170), .A(N5777), .B(N5776), .S0(N1135));
MXI2XL addgen2_A_I1511 (.Y(N1151), .A(N5868), .B(N5859), .S0(N4170));
MXI2XL addgen2_A_I1512 (.Y(N4179), .A(N5778), .B(N5777), .S0(N1135));
MXI2XL addgen2_A_I1513 (.Y(N1152), .A(N5868), .B(N5859), .S0(N4179));
MXI2XL addgen2_A_I1514 (.Y(N4188), .A(N5779), .B(N5778), .S0(N1135));
MXI2XL addgen2_A_I1515 (.Y(N1153), .A(N5868), .B(N5859), .S0(N4188));
MXI2XL addgen2_A_I1516 (.Y(N4197), .A(N5780), .B(N5779), .S0(N1135));
MXI2XL addgen2_A_I1517 (.Y(N1154), .A(N5868), .B(N5859), .S0(N4197));
MXI2XL addgen2_A_I1518 (.Y(N4206), .A(N5781), .B(N5780), .S0(N1135));
MXI2XL addgen2_A_I1519 (.Y(N1155), .A(N5868), .B(N5859), .S0(N4206));
MXI2XL addgen2_A_I1520 (.Y(N4215), .A(N5782), .B(N5781), .S0(N1135));
MXI2XL addgen2_A_I1521 (.Y(N1156), .A(N5868), .B(N5859), .S0(N4215));
MXI2XL addgen2_A_I1522 (.Y(N4224), .A(N5783), .B(N5782), .S0(N1135));
MXI2XL addgen2_A_I1523 (.Y(N1157), .A(N5868), .B(N5859), .S0(N4224));
MXI2XL addgen2_A_I1524 (.Y(N4233), .A(N5784), .B(N5783), .S0(N1135));
MXI2XL addgen2_A_I1525 (.Y(N1158), .A(N5868), .B(N5859), .S0(N4233));
MXI2XL addgen2_A_I1526 (.Y(N4242), .A(N5785), .B(N5784), .S0(N1135));
MXI2XL addgen2_A_I1527 (.Y(N1159), .A(N5868), .B(N5859), .S0(N4242));
MXI2XL addgen2_A_I1528 (.Y(N4251), .A(N5786), .B(N5785), .S0(N1135));
MXI2XL addgen2_A_I1529 (.Y(N1160), .A(N5868), .B(N5859), .S0(N4251));
MXI2XL addgen2_A_I1530 (.Y(N4260), .A(N5787), .B(N5786), .S0(N1135));
MXI2XL addgen2_A_I1531 (.Y(N1161), .A(N5868), .B(N5859), .S0(N4260));
MXI2XL addgen2_A_I1532 (.Y(N4269), .A(N5788), .B(N5787), .S0(N1135));
MXI2XL addgen2_A_I1533 (.Y(N1162), .A(N5868), .B(N5859), .S0(N4269));
NOR2BX1 addgen2_A_I1534 (.Y(N4278), .AN(N1135), .B(N5788));
MXI2XL addgen2_A_I1535 (.Y(N1163), .A(N5868), .B(N5859), .S0(N4278));
CLKINVX1 inst_cellmath__203_0_I2071 (.Y(N5869), .A(inst_cellmath__203_0_in0[7]));
INVXL inst_cellmath__203_0_I2072 (.Y(N5870), .A(N5869));
XNOR2X1 enc2_A_I1536 (.Y(N1167), .A(N5870), .B(N5844));
NAND2XL enc2_A_I1537 (.Y(N4287), .A(N5870), .B(N5844));
NOR2XL enc2_A_I1538 (.Y(N4289), .A(N5870), .B(N5844));
CLKINVX1 inst_cellmath__203_0_I2073 (.Y(N5871), .A(inst_cellmath__203_0_in0[8]));
INVXL inst_cellmath__203_0_I2074 (.Y(N5872), .A(N5871));
AND2XL enc2_A_I1539 (.Y(N1169), .A(N4287), .B(N5872));
OR2XL inst_cellmath__203_0_I2228 (.Y(N5887), .A(N4289), .B(N5872));
INVXL inst_cellmath__203_0_I2098 (.Y(N5896), .A(N1169));
NOR2XL addgen2_A_I1541 (.Y(N4300), .A(N5767), .B(N1167));
MXI2XL addgen2_A_I1542 (.Y(N1173), .A(N5896), .B(N5887), .S0(N4300));
MXI2XL addgen2_A_I1543 (.Y(N4309), .A(N5768), .B(N5767), .S0(N1167));
MXI2XL addgen2_A_I1544 (.Y(N1174), .A(N5896), .B(N5887), .S0(N4309));
MXI2XL addgen2_A_I1545 (.Y(N4318), .A(N5769), .B(N5768), .S0(N1167));
MXI2XL addgen2_A_I1546 (.Y(N1175), .A(N5896), .B(N5887), .S0(N4318));
MXI2XL addgen2_A_I1547 (.Y(N4327), .A(N5770), .B(N5769), .S0(N1167));
MXI2XL addgen2_A_I1548 (.Y(N1176), .A(N5896), .B(N5887), .S0(N4327));
MXI2XL addgen2_A_I1549 (.Y(N4336), .A(N5771), .B(N5770), .S0(N1167));
MXI2XL addgen2_A_I1550 (.Y(N1177), .A(N5896), .B(N5887), .S0(N4336));
MXI2XL addgen2_A_I1551 (.Y(N4345), .A(N5772), .B(N5771), .S0(N1167));
MXI2XL addgen2_A_I1552 (.Y(N1178), .A(N5896), .B(N5887), .S0(N4345));
MXI2XL addgen2_A_I1553 (.Y(N4354), .A(N5773), .B(N5772), .S0(N1167));
MXI2XL addgen2_A_I1554 (.Y(N1179), .A(N5896), .B(N5887), .S0(N4354));
MXI2XL addgen2_A_I1555 (.Y(N4363), .A(N5774), .B(N5773), .S0(N1167));
MXI2XL addgen2_A_I1556 (.Y(N1180), .A(N5896), .B(N5887), .S0(N4363));
MXI2XL addgen2_A_I1557 (.Y(N4372), .A(N5775), .B(N5774), .S0(N1167));
MXI2XL addgen2_A_I1558 (.Y(N1181), .A(N5896), .B(N5887), .S0(N4372));
MXI2XL addgen2_A_I1559 (.Y(N4381), .A(N5776), .B(N5775), .S0(N1167));
MXI2XL addgen2_A_I1560 (.Y(N1182), .A(N5896), .B(N5887), .S0(N4381));
MXI2XL addgen2_A_I1561 (.Y(N4390), .A(N5777), .B(N5776), .S0(N1167));
MXI2XL addgen2_A_I1562 (.Y(N1183), .A(N5896), .B(N5887), .S0(N4390));
MXI2XL addgen2_A_I1563 (.Y(N4399), .A(N5778), .B(N5777), .S0(N1167));
MXI2XL addgen2_A_I1564 (.Y(N1184), .A(N5896), .B(N5887), .S0(N4399));
MXI2XL addgen2_A_I1565 (.Y(N4408), .A(N5779), .B(N5778), .S0(N1167));
MXI2XL addgen2_A_I1566 (.Y(N1185), .A(N5896), .B(N5887), .S0(N4408));
MXI2XL addgen2_A_I1567 (.Y(N4417), .A(N5780), .B(N5779), .S0(N1167));
MXI2XL addgen2_A_I1568 (.Y(N1186), .A(N5896), .B(N5887), .S0(N4417));
MXI2XL addgen2_A_I1569 (.Y(N4426), .A(N5781), .B(N5780), .S0(N1167));
MXI2XL addgen2_A_I1570 (.Y(N1187), .A(N5896), .B(N5887), .S0(N4426));
MXI2XL addgen2_A_I1571 (.Y(N4435), .A(N5782), .B(N5781), .S0(N1167));
MXI2XL addgen2_A_I1572 (.Y(N1188), .A(N5896), .B(N5887), .S0(N4435));
MXI2XL addgen2_A_I1573 (.Y(N4444), .A(N5783), .B(N5782), .S0(N1167));
MXI2XL addgen2_A_I1574 (.Y(N1189), .A(N5896), .B(N5887), .S0(N4444));
MXI2XL addgen2_A_I1575 (.Y(N4453), .A(N5784), .B(N5783), .S0(N1167));
MXI2XL addgen2_A_I1576 (.Y(N1190), .A(N5896), .B(N5887), .S0(N4453));
MXI2XL addgen2_A_I1577 (.Y(N4462), .A(N5785), .B(N5784), .S0(N1167));
MXI2XL addgen2_A_I1578 (.Y(N1191), .A(N5896), .B(N5887), .S0(N4462));
MXI2XL addgen2_A_I1579 (.Y(N4471), .A(N5786), .B(N5785), .S0(N1167));
MXI2XL addgen2_A_I1580 (.Y(N1192), .A(N5896), .B(N5887), .S0(N4471));
MXI2XL addgen2_A_I1581 (.Y(N4480), .A(N5787), .B(N5786), .S0(N1167));
MXI2XL addgen2_A_I1582 (.Y(N1193), .A(N5896), .B(N5887), .S0(N4480));
MXI2XL addgen2_A_I1583 (.Y(N4489), .A(N5788), .B(N5787), .S0(N1167));
MXI2XL addgen2_A_I1584 (.Y(N1194), .A(N5896), .B(N5887), .S0(N4489));
NOR2BX1 addgen2_A_I1585 (.Y(N4498), .AN(N1167), .B(N5788));
MXI2XL addgen2_A_I1586 (.Y(N1195), .A(N5896), .B(N5887), .S0(N4498));
CLKINVX1 inst_cellmath__203_0_I2099 (.Y(N5897), .A(inst_cellmath__203_0_in0[9]));
INVXL inst_cellmath__203_0_I2100 (.Y(N5898), .A(N5897));
XNOR2X1 enc2_A_I1587 (.Y(N1199), .A(N5898), .B(N5872));
NAND2XL enc2_A_I1588 (.Y(N4507), .A(N5898), .B(N5872));
NOR2XL enc2_A_I1589 (.Y(N4509), .A(N5898), .B(N5872));
CLKINVX1 inst_cellmath__203_0_I2101 (.Y(N5899), .A(inst_cellmath__203_0_in0[10]));
INVXL inst_cellmath__203_0_I2102 (.Y(N5900), .A(N5899));
AND2XL enc2_A_I1590 (.Y(N1201), .A(N4507), .B(N5900));
OR2XL inst_cellmath__203_0_I2231 (.Y(N5915), .A(N4509), .B(N5900));
INVXL inst_cellmath__203_0_I2126 (.Y(N5924), .A(N1201));
NOR2XL addgen2_A_I1592 (.Y(N4520), .A(N5767), .B(N1199));
MXI2XL addgen2_A_I1593 (.Y(N1205), .A(N5924), .B(N5915), .S0(N4520));
MXI2XL addgen2_A_I1594 (.Y(N4529), .A(N5768), .B(N5767), .S0(N1199));
MXI2XL addgen2_A_I1595 (.Y(N1206), .A(N5924), .B(N5915), .S0(N4529));
MXI2XL addgen2_A_I1596 (.Y(N4538), .A(N5769), .B(N5768), .S0(N1199));
MXI2XL addgen2_A_I1597 (.Y(N1207), .A(N5924), .B(N5915), .S0(N4538));
MXI2XL addgen2_A_I1598 (.Y(N4547), .A(N5770), .B(N5769), .S0(N1199));
MXI2XL addgen2_A_I1599 (.Y(N1208), .A(N5924), .B(N5915), .S0(N4547));
MXI2XL addgen2_A_I1600 (.Y(N4556), .A(N5771), .B(N5770), .S0(N1199));
MXI2XL addgen2_A_I1601 (.Y(N1209), .A(N5924), .B(N5915), .S0(N4556));
MXI2XL addgen2_A_I1602 (.Y(N4565), .A(N5772), .B(N5771), .S0(N1199));
MXI2XL addgen2_A_I1603 (.Y(N1210), .A(N5924), .B(N5915), .S0(N4565));
MXI2XL addgen2_A_I1604 (.Y(N4574), .A(N5773), .B(N5772), .S0(N1199));
MXI2XL addgen2_A_I1605 (.Y(N1211), .A(N5924), .B(N5915), .S0(N4574));
MXI2XL addgen2_A_I1606 (.Y(N4583), .A(N5774), .B(N5773), .S0(N1199));
MXI2XL addgen2_A_I1607 (.Y(N1212), .A(N5924), .B(N5915), .S0(N4583));
MXI2XL addgen2_A_I1608 (.Y(N4592), .A(N5775), .B(N5774), .S0(N1199));
MXI2XL addgen2_A_I1609 (.Y(N1213), .A(N5924), .B(N5915), .S0(N4592));
MXI2XL addgen2_A_I1610 (.Y(N4601), .A(N5776), .B(N5775), .S0(N1199));
MXI2XL addgen2_A_I1611 (.Y(N1214), .A(N5924), .B(N5915), .S0(N4601));
MXI2XL addgen2_A_I1612 (.Y(N4610), .A(N5777), .B(N5776), .S0(N1199));
MXI2XL addgen2_A_I1613 (.Y(N1215), .A(N5924), .B(N5915), .S0(N4610));
MXI2XL addgen2_A_I1614 (.Y(N4619), .A(N5778), .B(N5777), .S0(N1199));
MXI2XL addgen2_A_I1615 (.Y(N1216), .A(N5924), .B(N5915), .S0(N4619));
MXI2XL addgen2_A_I1616 (.Y(N4628), .A(N5779), .B(N5778), .S0(N1199));
MXI2XL addgen2_A_I1617 (.Y(N1217), .A(N5924), .B(N5915), .S0(N4628));
MXI2XL addgen2_A_I1618 (.Y(N4637), .A(N5780), .B(N5779), .S0(N1199));
MXI2XL addgen2_A_I1619 (.Y(N1218), .A(N5924), .B(N5915), .S0(N4637));
MXI2XL addgen2_A_I1620 (.Y(N4646), .A(N5781), .B(N5780), .S0(N1199));
MXI2XL addgen2_A_I1621 (.Y(N1219), .A(N5924), .B(N5915), .S0(N4646));
MXI2XL addgen2_A_I1622 (.Y(N4655), .A(N5782), .B(N5781), .S0(N1199));
MXI2XL addgen2_A_I1623 (.Y(N1220), .A(N5924), .B(N5915), .S0(N4655));
MXI2XL addgen2_A_I1624 (.Y(N4664), .A(N5783), .B(N5782), .S0(N1199));
MXI2XL addgen2_A_I1625 (.Y(N1221), .A(N5924), .B(N5915), .S0(N4664));
MXI2XL addgen2_A_I1626 (.Y(N4673), .A(N5784), .B(N5783), .S0(N1199));
MXI2XL addgen2_A_I1627 (.Y(N1222), .A(N5924), .B(N5915), .S0(N4673));
MXI2XL addgen2_A_I1628 (.Y(N4682), .A(N5785), .B(N5784), .S0(N1199));
MXI2XL addgen2_A_I1629 (.Y(N1223), .A(N5924), .B(N5915), .S0(N4682));
MXI2XL addgen2_A_I1630 (.Y(N4691), .A(N5786), .B(N5785), .S0(N1199));
MXI2XL addgen2_A_I1631 (.Y(N1224), .A(N5924), .B(N5915), .S0(N4691));
MXI2XL addgen2_A_I1632 (.Y(N4700), .A(N5787), .B(N5786), .S0(N1199));
MXI2XL addgen2_A_I1633 (.Y(N1225), .A(N5924), .B(N5915), .S0(N4700));
MXI2XL addgen2_A_I1634 (.Y(N4709), .A(N5788), .B(N5787), .S0(N1199));
MXI2XL addgen2_A_I1635 (.Y(N1226), .A(N5924), .B(N5915), .S0(N4709));
NOR2BX1 addgen2_A_I1636 (.Y(N4718), .AN(N1199), .B(N5788));
MXI2XL addgen2_A_I1637 (.Y(N1227), .A(N5924), .B(N5915), .S0(N4718));
XNOR2X1 enc2_A_I1638 (.Y(N1231), .A(inst_cellmath__203_0_in0[11]), .B(N5900));
NAND2XL enc2_A_I1639 (.Y(N4727), .A(inst_cellmath__203_0_in0[11]), .B(N5900));
NOR2XL enc2_A_I1640 (.Y(N4729), .A(inst_cellmath__203_0_in0[11]), .B(N5900));
AND2XL enc2_A_I1641 (.Y(N1233), .A(N4727), .B(inst_cellmath__203_0_in0[12]));
OR2XL inst_cellmath__203_0_I2232 (.Y(N5939), .A(N4729), .B(inst_cellmath__203_0_in0[12]));
INVXL inst_cellmath__203_0_I2149 (.Y(N5947), .A(N1233));
NOR2XL addgen2_A_I1643 (.Y(N4740), .A(N5767), .B(N1231));
MXI2XL addgen2_A_I1644 (.Y(N1237), .A(N5947), .B(N5939), .S0(N4740));
MXI2XL addgen2_A_I1645 (.Y(N4749), .A(N5768), .B(N5767), .S0(N1231));
MXI2XL addgen2_A_I1646 (.Y(N1238), .A(N5947), .B(N5939), .S0(N4749));
MXI2XL addgen2_A_I1647 (.Y(N4758), .A(N5769), .B(N5768), .S0(N1231));
MXI2XL addgen2_A_I1648 (.Y(N1239), .A(N5947), .B(N5939), .S0(N4758));
MXI2XL addgen2_A_I1649 (.Y(N4767), .A(N5770), .B(N5769), .S0(N1231));
MXI2XL addgen2_A_I1650 (.Y(N1240), .A(N5947), .B(N5939), .S0(N4767));
MXI2XL addgen2_A_I1651 (.Y(N4776), .A(N5771), .B(N5770), .S0(N1231));
MXI2XL addgen2_A_I1652 (.Y(N1241), .A(N5947), .B(N5939), .S0(N4776));
MXI2XL addgen2_A_I1653 (.Y(N4785), .A(N5772), .B(N5771), .S0(N1231));
MXI2XL addgen2_A_I1654 (.Y(N1242), .A(N5947), .B(N5939), .S0(N4785));
MXI2XL addgen2_A_I1655 (.Y(N4794), .A(N5773), .B(N5772), .S0(N1231));
MXI2XL addgen2_A_I1656 (.Y(N1243), .A(N5947), .B(N5939), .S0(N4794));
MXI2XL addgen2_A_I1657 (.Y(N4803), .A(N5774), .B(N5773), .S0(N1231));
MXI2XL addgen2_A_I1658 (.Y(N1244), .A(N5947), .B(N5939), .S0(N4803));
MXI2XL addgen2_A_I1659 (.Y(N4812), .A(N5775), .B(N5774), .S0(N1231));
MXI2XL addgen2_A_I1660 (.Y(N1245), .A(N5947), .B(N5939), .S0(N4812));
MXI2XL addgen2_A_I1661 (.Y(N4821), .A(N5776), .B(N5775), .S0(N1231));
MXI2XL addgen2_A_I1662 (.Y(N1246), .A(N5947), .B(N5939), .S0(N4821));
MXI2XL addgen2_A_I1663 (.Y(N4830), .A(N5777), .B(N5776), .S0(N1231));
MXI2XL addgen2_A_I1664 (.Y(N1247), .A(N5947), .B(N5939), .S0(N4830));
MXI2XL addgen2_A_I1665 (.Y(N4839), .A(N5778), .B(N5777), .S0(N1231));
MXI2XL addgen2_A_I1666 (.Y(N1248), .A(N5947), .B(N5939), .S0(N4839));
MXI2XL addgen2_A_I1667 (.Y(N4848), .A(N5779), .B(N5778), .S0(N1231));
MXI2XL addgen2_A_I1668 (.Y(N1249), .A(N5947), .B(N5939), .S0(N4848));
MXI2XL addgen2_A_I1669 (.Y(N4857), .A(N5780), .B(N5779), .S0(N1231));
MXI2XL addgen2_A_I1670 (.Y(N1250), .A(N5947), .B(N5939), .S0(N4857));
MXI2XL addgen2_A_I1671 (.Y(N4866), .A(N5781), .B(N5780), .S0(N1231));
MXI2XL addgen2_A_I1672 (.Y(N1251), .A(N5947), .B(N5939), .S0(N4866));
MXI2XL addgen2_A_I1673 (.Y(N4875), .A(N5782), .B(N5781), .S0(N1231));
MXI2XL addgen2_A_I1674 (.Y(N1252), .A(N5947), .B(N5939), .S0(N4875));
MXI2XL addgen2_A_I1675 (.Y(N4884), .A(N5783), .B(N5782), .S0(N1231));
MXI2XL addgen2_A_I1676 (.Y(N1253), .A(N5947), .B(N5939), .S0(N4884));
MXI2XL addgen2_A_I1677 (.Y(N4893), .A(N5784), .B(N5783), .S0(N1231));
MXI2XL addgen2_A_I1678 (.Y(N1254), .A(N5947), .B(N5939), .S0(N4893));
MXI2XL addgen2_A_I1679 (.Y(N4902), .A(N5785), .B(N5784), .S0(N1231));
MXI2XL addgen2_A_I1680 (.Y(N1255), .A(N5947), .B(N5939), .S0(N4902));
MXI2XL addgen2_A_I1681 (.Y(N4911), .A(N5786), .B(N5785), .S0(N1231));
MXI2XL addgen2_A_I1682 (.Y(N1256), .A(N5947), .B(N5939), .S0(N4911));
MXI2XL addgen2_A_I1683 (.Y(N4920), .A(N5787), .B(N5786), .S0(N1231));
MXI2XL addgen2_A_I1684 (.Y(N1257), .A(N5947), .B(N5939), .S0(N4920));
MXI2XL addgen2_A_I1685 (.Y(N4929), .A(N5788), .B(N5787), .S0(N1231));
MXI2XL addgen2_A_I1686 (.Y(N1258), .A(N5947), .B(N5939), .S0(N4929));
NOR2BX1 addgen2_A_I1687 (.Y(N4938), .AN(N1231), .B(N5788));
MXI2XL addgen2_A_I1688 (.Y(N1259), .A(N5947), .B(N5939), .S0(N4938));
XNOR2X1 enc2_A_I1689 (.Y(N1263), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
NAND2XL enc2_A_I1690 (.Y(N4947), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
NOR2XL enc2_A_I1691 (.Y(N4949), .A(inst_cellmath__203_0_in0[13]), .B(inst_cellmath__203_0_in0[12]));
AND2XL enc2_A_I1692 (.Y(N1265), .A(N4947), .B(inst_cellmath__203_0_in0[14]));
OR2XL inst_cellmath__203_0_I2233 (.Y(N5962), .A(N4949), .B(inst_cellmath__203_0_in0[14]));
INVXL inst_cellmath__203_0_I2172 (.Y(N5970), .A(N1265));
NOR2XL addgen2_A_I1694 (.Y(N4960), .A(N5767), .B(N1263));
MXI2XL addgen2_A_I1695 (.Y(N1269), .A(N5970), .B(N5962), .S0(N4960));
MXI2XL addgen2_A_I1696 (.Y(N4969), .A(N5768), .B(N5767), .S0(N1263));
MXI2XL addgen2_A_I1697 (.Y(N1270), .A(N5970), .B(N5962), .S0(N4969));
MXI2XL addgen2_A_I1698 (.Y(N4978), .A(N5769), .B(N5768), .S0(N1263));
MXI2XL addgen2_A_I1699 (.Y(N1271), .A(N5970), .B(N5962), .S0(N4978));
MXI2XL addgen2_A_I1700 (.Y(N4987), .A(N5770), .B(N5769), .S0(N1263));
MXI2XL addgen2_A_I1701 (.Y(N1272), .A(N5970), .B(N5962), .S0(N4987));
MXI2XL addgen2_A_I1702 (.Y(N4996), .A(N5771), .B(N5770), .S0(N1263));
MXI2XL addgen2_A_I1703 (.Y(N1273), .A(N5970), .B(N5962), .S0(N4996));
MXI2XL addgen2_A_I1704 (.Y(N5005), .A(N5772), .B(N5771), .S0(N1263));
MXI2XL addgen2_A_I1705 (.Y(N1274), .A(N5970), .B(N5962), .S0(N5005));
MXI2XL addgen2_A_I1706 (.Y(N5014), .A(N5773), .B(N5772), .S0(N1263));
MXI2XL addgen2_A_I1707 (.Y(N1275), .A(N5970), .B(N5962), .S0(N5014));
MXI2XL addgen2_A_I1708 (.Y(N5023), .A(N5774), .B(N5773), .S0(N1263));
MXI2XL addgen2_A_I1709 (.Y(N1276), .A(N5970), .B(N5962), .S0(N5023));
MXI2XL addgen2_A_I1710 (.Y(N5032), .A(N5775), .B(N5774), .S0(N1263));
MXI2XL addgen2_A_I1711 (.Y(N1277), .A(N5970), .B(N5962), .S0(N5032));
MXI2XL addgen2_A_I1712 (.Y(N5041), .A(N5776), .B(N5775), .S0(N1263));
MXI2XL addgen2_A_I1713 (.Y(N1278), .A(N5970), .B(N5962), .S0(N5041));
MXI2XL addgen2_A_I1714 (.Y(N5050), .A(N5777), .B(N5776), .S0(N1263));
MXI2XL addgen2_A_I1715 (.Y(N1279), .A(N5970), .B(N5962), .S0(N5050));
MXI2XL addgen2_A_I1716 (.Y(N5059), .A(N5778), .B(N5777), .S0(N1263));
MXI2XL addgen2_A_I1717 (.Y(N1280), .A(N5970), .B(N5962), .S0(N5059));
MXI2XL addgen2_A_I1718 (.Y(N5068), .A(N5779), .B(N5778), .S0(N1263));
MXI2XL addgen2_A_I1719 (.Y(N1281), .A(N5970), .B(N5962), .S0(N5068));
MXI2XL addgen2_A_I1720 (.Y(N5077), .A(N5780), .B(N5779), .S0(N1263));
MXI2XL addgen2_A_I1721 (.Y(N1282), .A(N5970), .B(N5962), .S0(N5077));
MXI2XL addgen2_A_I1722 (.Y(N5086), .A(N5781), .B(N5780), .S0(N1263));
MXI2XL addgen2_A_I1723 (.Y(N1283), .A(N5970), .B(N5962), .S0(N5086));
MXI2XL addgen2_A_I1724 (.Y(N5095), .A(N5782), .B(N5781), .S0(N1263));
MXI2XL addgen2_A_I1725 (.Y(N1284), .A(N5970), .B(N5962), .S0(N5095));
MXI2XL addgen2_A_I1726 (.Y(N5104), .A(N5783), .B(N5782), .S0(N1263));
MXI2XL addgen2_A_I1727 (.Y(N1285), .A(N5970), .B(N5962), .S0(N5104));
MXI2XL addgen2_A_I1728 (.Y(N5113), .A(N5784), .B(N5783), .S0(N1263));
MXI2XL addgen2_A_I1729 (.Y(N1286), .A(N5970), .B(N5962), .S0(N5113));
MXI2XL addgen2_A_I1730 (.Y(N5122), .A(N5785), .B(N5784), .S0(N1263));
MXI2XL addgen2_A_I1731 (.Y(N1287), .A(N5970), .B(N5962), .S0(N5122));
MXI2XL addgen2_A_I1732 (.Y(N5131), .A(N5786), .B(N5785), .S0(N1263));
MXI2XL addgen2_A_I1733 (.Y(N1288), .A(N5970), .B(N5962), .S0(N5131));
MXI2XL addgen2_A_I1734 (.Y(N5140), .A(N5787), .B(N5786), .S0(N1263));
MXI2XL addgen2_A_I1735 (.Y(N1289), .A(N5970), .B(N5962), .S0(N5140));
MXI2XL addgen2_A_I1736 (.Y(N5149), .A(N5788), .B(N5787), .S0(N1263));
MXI2XL addgen2_A_I1737 (.Y(N1290), .A(N5970), .B(N5962), .S0(N5149));
NOR2BX1 addgen2_A_I1738 (.Y(N5158), .AN(N1263), .B(N5788));
MXI2XL addgen2_A_I1739 (.Y(N2112), .A(N5970), .B(N5962), .S0(N5158));
XNOR2X1 enc2_A_I1740 (.Y(N1295), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
NAND2XL enc2_A_I1741 (.Y(N5167), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
NOR2XL enc2_A_I1742 (.Y(N5169), .A(inst_cellmath__203_0_in0[15]), .B(inst_cellmath__203_0_in0[14]));
AND2XL enc2_A_I1743 (.Y(N1297), .A(N5167), .B(inst_cellmath__203_0_in4[0]));
OR2XL inst_cellmath__203_0_I2234 (.Y(N5985), .A(N5169), .B(inst_cellmath__203_0_in4[0]));
INVX2 inst_cellmath__203_0_I2195 (.Y(inst_cellmath__203_0_out1[42]), .A(N1297));
NOR2XL addgen2_A_I1745 (.Y(N5180), .A(N5767), .B(N1295));
MXI2XL addgen2_A_I1746 (.Y(N1301), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5180));
MXI2XL addgen2_A_I1747 (.Y(N5189), .A(N5768), .B(N5767), .S0(N1295));
MXI2XL addgen2_A_I1748 (.Y(N1302), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5189));
MXI2XL addgen2_A_I1749 (.Y(N5198), .A(N5769), .B(N5768), .S0(N1295));
MXI2XL addgen2_A_I1750 (.Y(N1303), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5198));
MXI2XL addgen2_A_I1751 (.Y(N5207), .A(N5770), .B(N5769), .S0(N1295));
MXI2XL addgen2_A_I1752 (.Y(N1304), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5207));
MXI2XL addgen2_A_I1753 (.Y(N5216), .A(N5771), .B(N5770), .S0(N1295));
MXI2XL addgen2_A_I1754 (.Y(N1305), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5216));
MXI2XL addgen2_A_I1755 (.Y(N5225), .A(N5772), .B(N5771), .S0(N1295));
MXI2XL addgen2_A_I1756 (.Y(N1306), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5225));
MXI2XL addgen2_A_I1757 (.Y(N5234), .A(N5773), .B(N5772), .S0(N1295));
MXI2XL addgen2_A_I1758 (.Y(N1307), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5234));
MXI2XL addgen2_A_I1759 (.Y(N5243), .A(N5774), .B(N5773), .S0(N1295));
MXI2XL addgen2_A_I1760 (.Y(N1308), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5243));
MXI2XL addgen2_A_I1761 (.Y(N5252), .A(N5775), .B(N5774), .S0(N1295));
MXI2XL addgen2_A_I1762 (.Y(N1309), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5252));
MXI2XL addgen2_A_I1763 (.Y(N5261), .A(N5776), .B(N5775), .S0(N1295));
MXI2XL addgen2_A_I1764 (.Y(N1310), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5261));
MXI2XL addgen2_A_I1765 (.Y(N5270), .A(N5777), .B(N5776), .S0(N1295));
MXI2XL addgen2_A_I1766 (.Y(N1311), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5270));
MXI2XL addgen2_A_I1767 (.Y(N5279), .A(N5778), .B(N5777), .S0(N1295));
MXI2XL addgen2_A_I1768 (.Y(N1312), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5279));
MXI2XL addgen2_A_I1769 (.Y(N5288), .A(N5779), .B(N5778), .S0(N1295));
MXI2XL addgen2_A_I1770 (.Y(N1313), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5288));
MXI2XL addgen2_A_I1771 (.Y(N5297), .A(N5780), .B(N5779), .S0(N1295));
MXI2XL addgen2_A_I1772 (.Y(N1314), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5297));
MXI2XL addgen2_A_I1773 (.Y(N5306), .A(N5781), .B(N5780), .S0(N1295));
MXI2XL addgen2_A_I1774 (.Y(N1315), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5306));
MXI2XL addgen2_A_I1775 (.Y(N5315), .A(N5782), .B(N5781), .S0(N1295));
MXI2XL addgen2_A_I1776 (.Y(N1316), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5315));
MXI2XL addgen2_A_I1777 (.Y(N5324), .A(N5783), .B(N5782), .S0(N1295));
MXI2XL addgen2_A_I1778 (.Y(N1317), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5324));
MXI2XL addgen2_A_I1779 (.Y(N5333), .A(N5784), .B(N5783), .S0(N1295));
MXI2XL addgen2_A_I1780 (.Y(N1318), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5333));
MXI2XL addgen2_A_I1781 (.Y(N5342), .A(N5785), .B(N5784), .S0(N1295));
MXI2XL addgen2_A_I1782 (.Y(N1319), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5342));
MXI2XL addgen2_A_I1783 (.Y(N5351), .A(N5786), .B(N5785), .S0(N1295));
MXI2XL addgen2_A_I1784 (.Y(N1320), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5351));
MXI2XL addgen2_A_I1785 (.Y(N5360), .A(N5787), .B(N5786), .S0(N1295));
MXI2XL addgen2_A_I1786 (.Y(N1321), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5360));
MXI2XL addgen2_A_I1787 (.Y(N5369), .A(N5788), .B(N5787), .S0(N1295));
MXI2XL addgen2_A_I1788 (.Y(N1322), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5369));
NOR2BX1 addgen2_A_I1789 (.Y(N5378), .AN(N1295), .B(N5788));
MXI2XL addgen2_A_I1790 (.Y(inst_cellmath__203_0_out0[42]), .A(inst_cellmath__203_0_out1[42]), .B(N5985), .S0(N5378));
ADDHX1 inst_cellmath__203_0_I684 (.CO(N1376), .S(inst_cellmath__203_0_out0[1]), .A(N518), .B(inst_cellmath__203_0_in1[19]));
ADDHX1 inst_cellmath__203_0_I685 (.CO(inst_cellmath__203_0_out1[3]), .S(inst_cellmath__203_0_out0[2]), .A(N520), .B(N1376));
ADDHX1 inst_cellmath__203_0_I686 (.CO(N1380), .S(N1379), .A(N522), .B(N591));
ADDFX1 inst_cellmath__203_0_I687 (.CO(N1382), .S(inst_cellmath__203_0_out0[3]), .A(N1379), .B(N567), .CI(N595));
ADDFX1 inst_cellmath__203_0_I688 (.CO(N1384), .S(inst_cellmath__203_0_out1[4]), .A(N524), .B(N1025), .CI(N568));
ADDFXL inst_cellmath__203_0_I689 (.CO(inst_cellmath__203_0_out1[5]), .S(inst_cellmath__203_0_out0[4]), .A(N596), .B(N1380), .CI(N1382));
ADDFX1 inst_cellmath__203_0_I690 (.CO(N1388), .S(N1387), .A(N1027), .B(inst_cellmath__203_0_in0[2]), .CI(N1077));
ADDFX1 inst_cellmath__203_0_I691 (.CO(N1390), .S(N1389), .A(N526), .B(N1387), .CI(N621));
ADDFXL inst_cellmath__203_0_I692 (.CO(N1392), .S(N1391), .A(N625), .B(N569), .CI(N597));
ADDFXL inst_cellmath__203_0_I693 (.CO(inst_cellmath__203_0_out1[6]), .S(inst_cellmath__203_0_out0[5]), .A(N1384), .B(N1389), .CI(N1391));
ADDFX1 inst_cellmath__203_0_I694 (.CO(N1396), .S(N1395), .A(N1078), .B(N1029), .CI(N1388));
ADDFX1 inst_cellmath__203_0_I695 (.CO(N1398), .S(N1397), .A(N528), .B(N1395), .CI(N570));
ADDFXL inst_cellmath__203_0_I696 (.CO(N1400), .S(N1399), .A(N1390), .B(N598), .CI(N626));
ADDFX1 inst_cellmath__203_0_I697 (.CO(inst_cellmath__203_0_out1[7]), .S(inst_cellmath__203_0_out0[6]), .A(N1392), .B(N1397), .CI(N1399));
ADDFX1 inst_cellmath__203_0_I698 (.CO(N1404), .S(N1403), .A(N1031), .B(N1105), .CI(N1079));
ADDFX1 inst_cellmath__203_0_I699 (.CO(N1406), .S(N1405), .A(N1403), .B(N1109), .CI(N1396));
ADDFX1 inst_cellmath__203_0_I700 (.CO(N1408), .S(N1407), .A(N1405), .B(N530), .CI(N651));
ADDFX1 inst_cellmath__203_0_I701 (.CO(N1410), .S(N1409), .A(N599), .B(N571), .CI(N655));
ADDFX1 inst_cellmath__203_0_I702 (.CO(N1412), .S(N1411), .A(N1407), .B(N627), .CI(N1398));
ADDFXL inst_cellmath__203_0_I703 (.CO(inst_cellmath__203_0_out1[8]), .S(inst_cellmath__203_0_out0[7]), .A(N1409), .B(N1400), .CI(N1411));
ADDFX1 inst_cellmath__203_0_I704 (.CO(N1416), .S(N1415), .A(N1080), .B(N1033), .CI(N1110));
ADDFX1 inst_cellmath__203_0_I705 (.CO(N1418), .S(N1417), .A(N1415), .B(N1404), .CI(N1406));
ADDFX1 inst_cellmath__203_0_I706 (.CO(N1420), .S(N1419), .A(N1417), .B(N532), .CI(N572));
ADDFX1 inst_cellmath__203_0_I707 (.CO(N1422), .S(N1421), .A(N1408), .B(N600), .CI(N656));
ADDFXL inst_cellmath__203_0_I708 (.CO(N1424), .S(N1423), .A(N1419), .B(N628), .CI(N1410));
ADDFXL inst_cellmath__203_0_I709 (.CO(inst_cellmath__203_0_out1[9]), .S(inst_cellmath__203_0_out0[8]), .A(N1421), .B(N1412), .CI(N1423));
ADDFX1 inst_cellmath__203_0_I710 (.CO(N1428), .S(N1427), .A(N1035), .B(N1137), .CI(N1111));
ADDFX1 inst_cellmath__203_0_I711 (.CO(N1430), .S(N1429), .A(N1141), .B(N1081), .CI(N1416));
ADDFX1 inst_cellmath__203_0_I712 (.CO(N1432), .S(N1431), .A(N1429), .B(N1427), .CI(N534));
ADDFX1 inst_cellmath__203_0_I713 (.CO(N1434), .S(N1433), .A(N681), .B(N1418), .CI(N1431));
ADDFX1 inst_cellmath__203_0_I714 (.CO(N1436), .S(N1435), .A(N601), .B(N573), .CI(N685));
ADDFX1 inst_cellmath__203_0_I715 (.CO(N1438), .S(N1437), .A(N629), .B(N657), .CI(N1433));
ADDFX1 inst_cellmath__203_0_I716 (.CO(N1440), .S(N1439), .A(N1422), .B(N1420), .CI(N1435));
ADDFXL inst_cellmath__203_0_I717 (.CO(inst_cellmath__203_0_out1[10]), .S(inst_cellmath__203_0_out0[9]), .A(N1424), .B(N1437), .CI(N1439));
ADDFX1 inst_cellmath__203_0_I718 (.CO(N1444), .S(N1443), .A(N1112), .B(N1037), .CI(N1142));
ADDFX1 inst_cellmath__203_0_I719 (.CO(N1446), .S(N1445), .A(N1428), .B(N1082), .CI(N1443));
ADDFX1 inst_cellmath__203_0_I720 (.CO(N1448), .S(N1447), .A(N1445), .B(N1430), .CI(N536));
ADDFX1 inst_cellmath__203_0_I721 (.CO(N1450), .S(N1449), .A(N1447), .B(N1432), .CI(N574));
ADDFX1 inst_cellmath__203_0_I722 (.CO(N1452), .S(N1451), .A(N686), .B(N602), .CI(N1434));
ADDFX1 inst_cellmath__203_0_I723 (.CO(N1454), .S(N1453), .A(N630), .B(N658), .CI(N1449));
ADDFXL inst_cellmath__203_0_I724 (.CO(N1456), .S(N1455), .A(N1438), .B(N1436), .CI(N1451));
ADDFXL inst_cellmath__203_0_I725 (.CO(inst_cellmath__203_0_out1[11]), .S(inst_cellmath__203_0_out0[10]), .A(N1440), .B(N1453), .CI(N1455));
ADDFX1 inst_cellmath__203_0_I726 (.CO(N1460), .S(N1459), .A(N1039), .B(N1169), .CI(N1083));
ADDFX1 inst_cellmath__203_0_I727 (.CO(N1462), .S(N1461), .A(N1113), .B(N1143), .CI(N1173));
ADDFX1 inst_cellmath__203_0_I728 (.CO(N1464), .S(N1463), .A(N1459), .B(N1444), .CI(N1461));
ADDFX1 inst_cellmath__203_0_I729 (.CO(N1466), .S(N1465), .A(N1463), .B(N1446), .CI(N538));
ADDFX1 inst_cellmath__203_0_I730 (.CO(N1468), .S(N1467), .A(N1465), .B(N1448), .CI(N711));
ADDFX1 inst_cellmath__203_0_I731 (.CO(N1470), .S(N1469), .A(N603), .B(N575), .CI(N687));
ADDFX1 inst_cellmath__203_0_I732 (.CO(N1472), .S(N1471), .A(N631), .B(N659), .CI(N715));
ADDFX1 inst_cellmath__203_0_I733 (.CO(N1474), .S(N1473), .A(N1450), .B(N1467), .CI(N1452));
ADDFX1 inst_cellmath__203_0_I734 (.CO(N1476), .S(N1475), .A(N1454), .B(N1469), .CI(N1471));
ADDFX1 inst_cellmath__203_0_I735 (.CO(inst_cellmath__203_0_out1[12]), .S(inst_cellmath__203_0_out0[11]), .A(N1456), .B(N1473), .CI(N1475));
ADDFX1 inst_cellmath__203_0_I736 (.CO(N1480), .S(N1479), .A(N1084), .B(N1041), .CI(N1144));
ADDFX1 inst_cellmath__203_0_I737 (.CO(N1482), .S(N1481), .A(N1174), .B(N1114), .CI(N1460));
ADDFX1 inst_cellmath__203_0_I738 (.CO(N1484), .S(N1483), .A(N1479), .B(N1462), .CI(N1481));
ADDFX1 inst_cellmath__203_0_I739 (.CO(N1486), .S(N1485), .A(N540), .B(N1464), .CI(N1483));
ADDFX1 inst_cellmath__203_0_I740 (.CO(N1488), .S(N1487), .A(N576), .B(N1466), .CI(N1485));
ADDFX1 inst_cellmath__203_0_I741 (.CO(N1490), .S(N1489), .A(N688), .B(N604), .CI(N1468));
ADDFX1 inst_cellmath__203_0_I742 (.CO(N1492), .S(N1491), .A(N632), .B(N660), .CI(N716));
ADDFX1 inst_cellmath__203_0_I743 (.CO(N1494), .S(N1493), .A(N1487), .B(N1470), .CI(N1472));
ADDFX1 inst_cellmath__203_0_I744 (.CO(N1496), .S(N1495), .A(N1491), .B(N1489), .CI(N1474));
ADDFX1 inst_cellmath__203_0_I745 (.CO(inst_cellmath__203_0_out1[13]), .S(inst_cellmath__203_0_out0[12]), .A(N1476), .B(N1493), .CI(N1495));
ADDFX1 inst_cellmath__203_0_I746 (.CO(N1500), .S(N1499), .A(N1043), .B(N1201), .CI(N1115));
ADDFX1 inst_cellmath__203_0_I747 (.CO(N1502), .S(N1501), .A(N1145), .B(N1175), .CI(N1205));
ADDFX1 inst_cellmath__203_0_I748 (.CO(N1504), .S(N1503), .A(N1480), .B(N1085), .CI(N1499));
ADDFXL inst_cellmath__203_0_I749 (.CO(N1506), .S(N1505), .A(N1482), .B(N1501), .CI(N1503));
ADDFX1 inst_cellmath__203_0_I750 (.CO(N1508), .S(N1507), .A(N1484), .B(N542), .CI(N1505));
ADDFX1 inst_cellmath__203_0_I751 (.CO(N1510), .S(N1509), .A(N577), .B(N1486), .CI(N741));
ADDFX1 inst_cellmath__203_0_I752 (.CO(N1512), .S(N1511), .A(N1507), .B(N605), .CI(N689));
ADDFX1 inst_cellmath__203_0_I753 (.CO(N1514), .S(N1513), .A(N633), .B(N661), .CI(N717));
ADDFX1 inst_cellmath__203_0_I754 (.CO(N1516), .S(N1515), .A(N1488), .B(N745), .CI(N1509));
ADDFX1 inst_cellmath__203_0_I755 (.CO(N1518), .S(N1517), .A(N1492), .B(N1490), .CI(N1511));
ADDFXL inst_cellmath__203_0_I756 (.CO(N1520), .S(N1519), .A(N1494), .B(N1513), .CI(N1515));
ADDFX1 inst_cellmath__203_0_I757 (.CO(inst_cellmath__203_0_out1[14]), .S(inst_cellmath__203_0_out0[13]), .A(N1496), .B(N1517), .CI(N1519));
ADDFX1 inst_cellmath__203_0_I758 (.CO(N1524), .S(N1523), .A(N1116), .B(N1045), .CI(N1176));
ADDFX1 inst_cellmath__203_0_I759 (.CO(N1526), .S(N1525), .A(N1206), .B(N1146), .CI(N1086));
ADDFXL inst_cellmath__203_0_I760 (.CO(N1528), .S(N1527), .A(N1502), .B(N1500), .CI(N1523));
ADDFXL inst_cellmath__203_0_I761 (.CO(N1530), .S(N1529), .A(N1504), .B(N1525), .CI(N1527));
ADDFX1 inst_cellmath__203_0_I762 (.CO(N1532), .S(N1531), .A(N1506), .B(N544), .CI(N1529));
ADDFXL inst_cellmath__203_0_I763 (.CO(N1534), .S(N1533), .A(N1508), .B(N578), .CI(N606));
ADDFX1 inst_cellmath__203_0_I764 (.CO(N1536), .S(N1535), .A(N662), .B(N690), .CI(N634));
ADDFX1 inst_cellmath__203_0_I765 (.CO(N1538), .S(N1537), .A(N718), .B(N1531), .CI(N746));
ADDFXL inst_cellmath__203_0_I766 (.CO(N1540), .S(N1539), .A(N1512), .B(N1510), .CI(N1533));
ADDFXL inst_cellmath__203_0_I767 (.CO(N1542), .S(N1541), .A(N1535), .B(N1514), .CI(N1516));
ADDFX1 inst_cellmath__203_0_I768 (.CO(N1544), .S(N1543), .A(N1518), .B(N1537), .CI(N1539));
ADDFXL inst_cellmath__203_0_I769 (.CO(inst_cellmath__203_0_out1[15]), .S(inst_cellmath__203_0_out0[14]), .A(N1541), .B(N1520), .CI(N1543));
ADDHX1 inst_cellmath__203_0_I770 (.CO(N1548), .S(N1547), .A(N1233), .B(N1047));
ADDFX1 inst_cellmath__203_0_I771 (.CO(N1550), .S(N1549), .A(N1147), .B(N1547), .CI(N1087));
ADDFX1 inst_cellmath__203_0_I772 (.CO(N1552), .S(N1551), .A(N1177), .B(N1207), .CI(N1237));
ADDFX1 inst_cellmath__203_0_I773 (.CO(N1554), .S(N1553), .A(N1524), .B(N1117), .CI(N1526));
ADDFX1 inst_cellmath__203_0_I774 (.CO(N1556), .S(N1555), .A(N1551), .B(N1549), .CI(N1528));
ADDFXL inst_cellmath__203_0_I775 (.CO(N1558), .S(N1557), .A(N546), .B(N1553), .CI(N1530));
ADDFX1 inst_cellmath__203_0_I776 (.CO(N1560), .S(N1559), .A(N579), .B(N1555), .CI(N779));
ADDFXL inst_cellmath__203_0_I777 (.CO(N1562), .S(N1561), .A(N1557), .B(N1532), .CI(N607));
ADDFX1 inst_cellmath__203_0_I778 (.CO(N1564), .S(N1563), .A(N663), .B(N691), .CI(N635));
ADDFX1 inst_cellmath__203_0_I779 (.CO(N1566), .S(N1565), .A(N747), .B(N719), .CI(N1534));
ADDFXL inst_cellmath__203_0_I780 (.CO(N1568), .S(N1567), .A(N1536), .B(N1559), .CI(N1561));
ADDFXL inst_cellmath__203_0_I781 (.CO(N1570), .S(N1569), .A(N1563), .B(N1538), .CI(N1540));
ADDFXL inst_cellmath__203_0_I782 (.CO(N1572), .S(N1571), .A(N1567), .B(N1565), .CI(N1542));
ADDFXL inst_cellmath__203_0_I783 (.CO(inst_cellmath__203_0_out1[16]), .S(inst_cellmath__203_0_out0[15]), .A(N1544), .B(N1569), .CI(N1571));
ADDFX1 inst_cellmath__203_0_I784 (.CO(N1576), .S(N1575), .A(N1548), .B(N1049), .CI(N1148));
ADDFX1 inst_cellmath__203_0_I785 (.CO(N1578), .S(N1577), .A(N1208), .B(N1088), .CI(N1118));
ADDFX1 inst_cellmath__203_0_I786 (.CO(N1580), .S(N1579), .A(N1238), .B(N1178), .CI(N1550));
ADDFX1 inst_cellmath__203_0_I787 (.CO(N1582), .S(N1581), .A(N1575), .B(N1552), .CI(N1577));
ADDFXL inst_cellmath__203_0_I788 (.CO(N1584), .S(N1583), .A(N1579), .B(N1554), .CI(N1581));
ADDFXL inst_cellmath__203_0_I789 (.CO(N1586), .S(N1585), .A(N1556), .B(N548), .CI(N1583));
ADDFXL inst_cellmath__203_0_I790 (.CO(N1588), .S(N1587), .A(N580), .B(N1558), .CI(N608));
ADDFXL inst_cellmath__203_0_I791 (.CO(N1590), .S(N1589), .A(N692), .B(N781), .CI(N664));
ADDFXL inst_cellmath__203_0_I792 (.CO(N1592), .S(N1591), .A(N1585), .B(N636), .CI(N720));
ADDFX1 inst_cellmath__203_0_I793 (.CO(N1594), .S(N1593), .A(N1560), .B(N748), .CI(N1562));
ADDFXL inst_cellmath__203_0_I794 (.CO(N1596), .S(N1595), .A(N1587), .B(N1564), .CI(N1589));
ADDFXL inst_cellmath__203_0_I795 (.CO(N1598), .S(N1597), .A(N1566), .B(N1591), .CI(N1593));
ADDFXL inst_cellmath__203_0_I796 (.CO(N1600), .S(N1599), .A(N1595), .B(N1568), .CI(N1570));
ADDFXL inst_cellmath__203_0_I797 (.CO(inst_cellmath__203_0_out1[17]), .S(inst_cellmath__203_0_out0[16]), .A(N1572), .B(N1597), .CI(N1599));
ADDFX1 inst_cellmath__203_0_I798 (.CO(N1604), .S(N1603), .A(N1051), .B(N1265), .CI(N1089));
ADDFX1 inst_cellmath__203_0_I799 (.CO(N1606), .S(N1605), .A(N1239), .B(N1179), .CI(N1209));
ADDFX1 inst_cellmath__203_0_I800 (.CO(N1608), .S(N1607), .A(N1269), .B(N1119), .CI(N1149));
ADDFX1 inst_cellmath__203_0_I801 (.CO(N1610), .S(N1609), .A(N1578), .B(N1576), .CI(N1603));
ADDFX1 inst_cellmath__203_0_I802 (.CO(N1612), .S(N1611), .A(N1607), .B(N1605), .CI(N1580));
ADDFXL inst_cellmath__203_0_I803 (.CO(N1614), .S(N1613), .A(N1609), .B(N1582), .CI(N550));
ADDFX1 inst_cellmath__203_0_I804 (.CO(N1616), .S(N1615), .A(N1584), .B(N1611), .CI(N1613));
ADDFXL inst_cellmath__203_0_I805 (.CO(N1618), .S(N1617), .A(N1586), .B(N581), .CI(N609));
ADDFXL inst_cellmath__203_0_I806 (.CO(N1620), .S(N1619), .A(N693), .B(N783), .CI(N665));
ADDFX1 inst_cellmath__203_0_I807 (.CO(N1622), .S(N1621), .A(N721), .B(N637), .CI(N1615));
ADDFX1 inst_cellmath__203_0_I808 (.CO(N1624), .S(N1623), .A(N1588), .B(N749), .CI(N1590));
ADDFXL inst_cellmath__203_0_I809 (.CO(N1626), .S(N1625), .A(N1619), .B(N1592), .CI(N1617));
ADDFX1 inst_cellmath__203_0_I810 (.CO(N1628), .S(N1627), .A(N1621), .B(N1594), .CI(N1596));
ADDFXL inst_cellmath__203_0_I811 (.CO(N1630), .S(N1629), .A(N1625), .B(N1623), .CI(N1598));
ADDFXL inst_cellmath__203_0_I812 (.CO(inst_cellmath__203_0_out1[18]), .S(inst_cellmath__203_0_out0[17]), .A(N1600), .B(N1627), .CI(N1629));
ADDFX1 inst_cellmath__203_0_I813 (.CO(N1634), .S(N1633), .A(N1180), .B(N1053), .CI(N1210));
ADDFX1 inst_cellmath__203_0_I814 (.CO(N1636), .S(N1635), .A(N1240), .B(N1120), .CI(N1150));
ADDFXL inst_cellmath__203_0_I815 (.CO(N1638), .S(N1637), .A(N1270), .B(N1090), .CI(N1604));
ADDFX1 inst_cellmath__203_0_I816 (.CO(N1640), .S(N1639), .A(N1608), .B(N1606), .CI(N1633));
ADDFX1 inst_cellmath__203_0_I817 (.CO(N1642), .S(N1641), .A(N1637), .B(N1635), .CI(N1610));
ADDFXL inst_cellmath__203_0_I818 (.CO(N1644), .S(N1643), .A(N1639), .B(N1612), .CI(N552));
ADDFX1 inst_cellmath__203_0_I819 (.CO(N1646), .S(N1645), .A(N1614), .B(N1641), .CI(N1643));
ADDFXL inst_cellmath__203_0_I820 (.CO(N1648), .S(N1647), .A(N1616), .B(N582), .CI(N610));
ADDFXL inst_cellmath__203_0_I821 (.CO(N1650), .S(N1649), .A(N694), .B(N785), .CI(N666));
ADDFXL inst_cellmath__203_0_I822 (.CO(N1652), .S(N1651), .A(N722), .B(N638), .CI(N1645));
ADDFX1 inst_cellmath__203_0_I823 (.CO(N1654), .S(N1653), .A(N1618), .B(N750), .CI(N1620));
ADDFX1 inst_cellmath__203_0_I824 (.CO(N1656), .S(N1655), .A(N1647), .B(N1622), .CI(N1649));
ADDFXL inst_cellmath__203_0_I825 (.CO(N1658), .S(N1657), .A(N1624), .B(N1651), .CI(N1626));
ADDFX1 inst_cellmath__203_0_I826 (.CO(N1660), .S(N1659), .A(N1655), .B(N1653), .CI(N1628));
ADDFX1 inst_cellmath__203_0_I827 (.CO(inst_cellmath__203_0_out1[19]), .S(inst_cellmath__203_0_out0[18]), .A(N1630), .B(N1657), .CI(N1659));
ADDFX1 inst_cellmath__203_0_I828 (.CO(N1664), .S(N1663), .A(N1055), .B(N1297), .CI(N1121));
ADDFX1 inst_cellmath__203_0_I829 (.CO(N1666), .S(N1665), .A(N1271), .B(N1211), .CI(N1241));
ADDFX1 inst_cellmath__203_0_I830 (.CO(N1668), .S(N1667), .A(N1091), .B(N1151), .CI(N1181));
ADDFX1 inst_cellmath__203_0_I831 (.CO(N1670), .S(N1669), .A(N1634), .B(N1301), .CI(N1636));
ADDFXL inst_cellmath__203_0_I832 (.CO(N1672), .S(N1671), .A(N1665), .B(N1663), .CI(N1638));
ADDFX1 inst_cellmath__203_0_I833 (.CO(N1674), .S(N1673), .A(N1640), .B(N1667), .CI(N1669));
ADDFXL inst_cellmath__203_0_I834 (.CO(N1676), .S(N1675), .A(N1671), .B(N1642), .CI(N554));
ADDFXL inst_cellmath__203_0_I835 (.CO(N1678), .S(N1677), .A(N1644), .B(N1673), .CI(N1675));
ADDFXL inst_cellmath__203_0_I836 (.CO(N1680), .S(N1679), .A(N611), .B(N583), .CI(N1646));
ADDFXL inst_cellmath__203_0_I837 (.CO(N1682), .S(N1681), .A(N695), .B(N787), .CI(N667));
ADDFX1 inst_cellmath__203_0_I838 (.CO(N1684), .S(N1683), .A(N723), .B(N639), .CI(N1677));
ADDFX1 inst_cellmath__203_0_I839 (.CO(N1686), .S(N1685), .A(N1648), .B(N751), .CI(N1650));
ADDFXL inst_cellmath__203_0_I840 (.CO(N1688), .S(N1687), .A(N1679), .B(N1652), .CI(N1681));
ADDFXL inst_cellmath__203_0_I841 (.CO(N1690), .S(N1689), .A(N1654), .B(N1683), .CI(N1656));
ADDFXL inst_cellmath__203_0_I842 (.CO(N1692), .S(N1691), .A(N1687), .B(N1685), .CI(N1658));
ADDFXL inst_cellmath__203_0_I843 (.CO(inst_cellmath__203_0_out1[20]), .S(inst_cellmath__203_0_out0[19]), .A(N1660), .B(N1689), .CI(N1691));
INVXL fap1_A_I1791 (.Y(N5387), .A(N1698));
ADDFX1 fap1_A_I1792 (.CO(N1696), .S(N1695), .A(N1152), .B(N1212), .CI(N5387));
ADDFX1 inst_cellmath__203_0_I845 (.CO(N1700), .S(N1699), .A(N1242), .B(N1272), .CI(N1182));
ADDFX1 inst_cellmath__203_0_I846 (.CO(N1702), .S(N1701), .A(N1092), .B(N1122), .CI(N1302));
ADDFX1 inst_cellmath__203_0_I847 (.CO(N1704), .S(N1703), .A(N1666), .B(N1664), .CI(N1668));
ADDFX1 inst_cellmath__203_0_I848 (.CO(N1706), .S(N1705), .A(N1701), .B(N1699), .CI(N1695));
ADDFX1 inst_cellmath__203_0_I849 (.CO(N1708), .S(N1707), .A(N1672), .B(N1670), .CI(N1703));
ADDFX1 inst_cellmath__203_0_I850 (.CO(N1710), .S(N1709), .A(N1705), .B(N5650), .CI(N1674));
ADDFX1 inst_cellmath__203_0_I851 (.CO(N1712), .S(N1711), .A(N1676), .B(N1707), .CI(N1709));
ADDFXL inst_cellmath__203_0_I852 (.CO(N1714), .S(N1713), .A(N612), .B(N584), .CI(N696));
ADDFXL inst_cellmath__203_0_I853 (.CO(N1716), .S(N1715), .A(N1678), .B(N789), .CI(N668));
ADDFX1 inst_cellmath__203_0_I854 (.CO(N1718), .S(N1717), .A(N724), .B(N640), .CI(N752));
ADDFX1 inst_cellmath__203_0_I855 (.CO(N1720), .S(N1719), .A(N1680), .B(N1711), .CI(N1682));
ADDFXL inst_cellmath__203_0_I856 (.CO(N1722), .S(N1721), .A(N1713), .B(N1684), .CI(N1715));
ADDFXL inst_cellmath__203_0_I857 (.CO(N1724), .S(N1723), .A(N1717), .B(N1686), .CI(N1688));
ADDFXL inst_cellmath__203_0_I858 (.CO(N1726), .S(N1725), .A(N1721), .B(N1719), .CI(N1690));
ADDFXL inst_cellmath__203_0_I859 (.CO(inst_cellmath__203_0_out1[21]), .S(inst_cellmath__203_0_out0[20]), .A(N1692), .B(N1723), .CI(N1725));
INVXL fap1_A_I1793 (.Y(N5396), .A(N1732));
ADDFX1 fap1_A_I1794 (.CO(N1730), .S(N1729), .A(N1153), .B(N1698), .CI(N5396));
ADDFX1 inst_cellmath__203_0_I861 (.CO(N1734), .S(N1733), .A(N1093), .B(N1243), .CI(N1273));
ADDFX1 inst_cellmath__203_0_I862 (.CO(N1736), .S(N1735), .A(N1183), .B(N1303), .CI(N1123));
ADDFX1 inst_cellmath__203_0_I863 (.CO(N1738), .S(N1737), .A(N1696), .B(N1213), .CI(N1702));
ADDFX1 inst_cellmath__203_0_I864 (.CO(N1740), .S(N1739), .A(N1733), .B(N1700), .CI(N1735));
ADDFX1 inst_cellmath__203_0_I865 (.CO(N1742), .S(N1741), .A(N1704), .B(N1729), .CI(N1737));
ADDFX1 inst_cellmath__203_0_I866 (.CO(N1744), .S(N1743), .A(N1739), .B(N1706), .CI(N1708));
ADDFX1 inst_cellmath__203_0_I867 (.CO(N1746), .S(N1745), .A(N1710), .B(N1741), .CI(N585));
ADDFX1 inst_cellmath__203_0_I868 (.CO(N1748), .S(N1747), .A(N613), .B(N1743), .CI(N697));
ADDFX1 inst_cellmath__203_0_I869 (.CO(N1750), .S(N1749), .A(N669), .B(N791), .CI(N641));
ADDFX1 inst_cellmath__203_0_I870 (.CO(N1752), .S(N1751), .A(N725), .B(N1712), .CI(N753));
ADDFX1 inst_cellmath__203_0_I871 (.CO(N1754), .S(N1753), .A(N1714), .B(N1745), .CI(N1716));
ADDFXL inst_cellmath__203_0_I872 (.CO(N1756), .S(N1755), .A(N1718), .B(N1747), .CI(N1749));
ADDFXL inst_cellmath__203_0_I873 (.CO(N1758), .S(N1757), .A(N1751), .B(N1720), .CI(N1722));
ADDFXL inst_cellmath__203_0_I874 (.CO(N1760), .S(N1759), .A(N1755), .B(N1753), .CI(N1724));
ADDFXL inst_cellmath__203_0_I875 (.CO(inst_cellmath__203_0_out1[22]), .S(inst_cellmath__203_0_out0[21]), .A(N1726), .B(N1757), .CI(N1759));
ADDFX1 inst_cellmath__203_0_I876 (.CO(N1764), .S(N1763), .A(N1061), .B(N1732), .CI(N1094));
ADDFX1 inst_cellmath__203_0_I877 (.CO(N1766), .S(N1765), .A(N1184), .B(N1244), .CI(N1274));
ADDFX1 inst_cellmath__203_0_I878 (.CO(N1768), .S(N1767), .A(N1154), .B(N1304), .CI(N1214));
ADDFX1 inst_cellmath__203_0_I879 (.CO(N1770), .S(N1769), .A(N1730), .B(N1124), .CI(N1736));
ADDFX1 inst_cellmath__203_0_I880 (.CO(N1772), .S(N1771), .A(N1763), .B(N1734), .CI(N1765));
ADDFX1 inst_cellmath__203_0_I881 (.CO(N1774), .S(N1773), .A(N1738), .B(N1767), .CI(N1769));
ADDFX1 inst_cellmath__203_0_I882 (.CO(N1776), .S(N1775), .A(N1771), .B(N1740), .CI(N1742));
ADDFXL inst_cellmath__203_0_I883 (.CO(N1778), .S(N1777), .A(N5666), .B(N1773), .CI(N1744));
ADDFXL inst_cellmath__203_0_I884 (.CO(N1780), .S(N1779), .A(N614), .B(N1775), .CI(N698));
ADDFXL inst_cellmath__203_0_I885 (.CO(N1782), .S(N1781), .A(N670), .B(N793), .CI(N642));
ADDFX1 inst_cellmath__203_0_I886 (.CO(N1784), .S(N1783), .A(N1777), .B(N726), .CI(N1746));
ADDFXL inst_cellmath__203_0_I887 (.CO(N1786), .S(N1785), .A(N1748), .B(N754), .CI(N1750));
ADDFXL inst_cellmath__203_0_I888 (.CO(N1788), .S(N1787), .A(N1752), .B(N1779), .CI(N1781));
ADDFXL inst_cellmath__203_0_I889 (.CO(N1790), .S(N1789), .A(N1754), .B(N1783), .CI(N1785));
ADDFXL inst_cellmath__203_0_I890 (.CO(N1792), .S(N1791), .A(N1787), .B(N1756), .CI(N1758));
ADDFXL inst_cellmath__203_0_I891 (.CO(inst_cellmath__203_0_out1[23]), .S(inst_cellmath__203_0_out0[22]), .A(N1760), .B(N1789), .CI(N1791));
INVXL fap1_A_I1795 (.Y(N5405), .A(N1798));
ADDFX1 fap1_A_I1796 (.CO(N1796), .S(N1795), .A(N1095), .B(N1185), .CI(N5405));
ADDFX1 inst_cellmath__203_0_I893 (.CO(N1800), .S(N1799), .A(N1125), .B(N1275), .CI(N1305));
ADDFX1 inst_cellmath__203_0_I894 (.CO(N1802), .S(N1801), .A(N1155), .B(N1215), .CI(N1245));
ADDFX1 inst_cellmath__203_0_I895 (.CO(N1804), .S(N1803), .A(N1766), .B(N1764), .CI(N1768));
ADDFX1 inst_cellmath__203_0_I896 (.CO(N1806), .S(N1805), .A(N1795), .B(N1799), .CI(N1801));
ADDFX1 inst_cellmath__203_0_I897 (.CO(N1808), .S(N1807), .A(N1772), .B(N1770), .CI(N1803));
ADDFX1 inst_cellmath__203_0_I898 (.CO(N1810), .S(N1809), .A(N1774), .B(N1805), .CI(N1807));
ADDFXL inst_cellmath__203_0_I899 (.CO(N1812), .S(N1811), .A(N615), .B(N1776), .CI(N1778));
ADDFX1 inst_cellmath__203_0_I900 (.CO(N1814), .S(N1813), .A(N699), .B(N795), .CI(N1809));
ADDFX1 inst_cellmath__203_0_I901 (.CO(N1816), .S(N1815), .A(N643), .B(N671), .CI(N727));
ADDFXL inst_cellmath__203_0_I902 (.CO(N1818), .S(N1817), .A(N1780), .B(N755), .CI(N1782));
ADDFXL inst_cellmath__203_0_I903 (.CO(N1820), .S(N1819), .A(N1811), .B(N1784), .CI(N1813));
ADDFXL inst_cellmath__203_0_I904 (.CO(N1822), .S(N1821), .A(N1786), .B(N1815), .CI(N1817));
ADDFXL inst_cellmath__203_0_I905 (.CO(N1824), .S(N1823), .A(N1819), .B(N1788), .CI(N1790));
ADDFXL inst_cellmath__203_0_I906 (.CO(inst_cellmath__203_0_out1[24]), .S(inst_cellmath__203_0_out0[23]), .A(N1792), .B(N1821), .CI(N1823));
INVXL fap1_A_I1797 (.Y(N5414), .A(N1830));
ADDFX1 fap1_A_I1798 (.CO(N1828), .S(N1827), .A(N1096), .B(N1798), .CI(N5414));
ADDFX1 inst_cellmath__203_0_I908 (.CO(N1832), .S(N1831), .A(N1276), .B(N1126), .CI(N1306));
ADDFX1 inst_cellmath__203_0_I909 (.CO(N1834), .S(N1833), .A(N1186), .B(N1216), .CI(N1156));
ADDFX1 inst_cellmath__203_0_I910 (.CO(N1836), .S(N1835), .A(N1796), .B(N1246), .CI(N1800));
ADDFX1 inst_cellmath__203_0_I911 (.CO(N1838), .S(N1837), .A(N1831), .B(N1802), .CI(N1833));
ADDFX1 inst_cellmath__203_0_I912 (.CO(N1840), .S(N1839), .A(N1804), .B(N1827), .CI(N1835));
ADDFXL inst_cellmath__203_0_I913 (.CO(N1842), .S(N1841), .A(N1837), .B(N1806), .CI(N1808));
ADDFX1 inst_cellmath__203_0_I914 (.CO(N1844), .S(N1843), .A(N5683), .B(N1839), .CI(N1841));
ADDFX1 inst_cellmath__203_0_I915 (.CO(N1846), .S(N1845), .A(N797), .B(N1810), .CI(N700));
ADDFX1 inst_cellmath__203_0_I916 (.CO(N1848), .S(N1847), .A(N644), .B(N672), .CI(N728));
ADDFXL inst_cellmath__203_0_I917 (.CO(N1850), .S(N1849), .A(N1843), .B(N756), .CI(N1812));
ADDFX1 inst_cellmath__203_0_I918 (.CO(N1852), .S(N1851), .A(N1816), .B(N1814), .CI(N1845));
ADDFX1 inst_cellmath__203_0_I919 (.CO(N1854), .S(N1853), .A(N1818), .B(N1847), .CI(N1849));
ADDFXL inst_cellmath__203_0_I920 (.CO(N1856), .S(N1855), .A(N1851), .B(N1820), .CI(N1822));
ADDFXL inst_cellmath__203_0_I921 (.CO(inst_cellmath__203_0_out1[25]), .S(inst_cellmath__203_0_out0[24]), .A(N1824), .B(N1853), .CI(N1855));
XNOR2X1 hap1_A_I1799 (.Y(N1859), .A(N1067), .B(N1830));
OR2XL hap1_A_I1800 (.Y(N1860), .A(N1067), .B(N1830));
ADDFX1 inst_cellmath__203_0_I923 (.CO(N1864), .S(N1863), .A(N1217), .B(N1859), .CI(N1307));
ADDFX1 inst_cellmath__203_0_I924 (.CO(N1866), .S(N1865), .A(N1127), .B(N1097), .CI(N1157));
ADDFX1 inst_cellmath__203_0_I925 (.CO(N1868), .S(N1867), .A(N1187), .B(N1247), .CI(N1277));
ADDFX1 inst_cellmath__203_0_I926 (.CO(N1870), .S(N1869), .A(N1832), .B(N1828), .CI(N1834));
ADDFX1 inst_cellmath__203_0_I927 (.CO(N1872), .S(N1871), .A(N1865), .B(N1863), .CI(N1867));
ADDFX1 inst_cellmath__203_0_I928 (.CO(N1874), .S(N1873), .A(N1869), .B(N1836), .CI(N1838));
ADDFX1 inst_cellmath__203_0_I929 (.CO(N1876), .S(N1875), .A(N1840), .B(N1871), .CI(N1873));
ADDFX1 inst_cellmath__203_0_I930 (.CO(N1878), .S(N1877), .A(N799), .B(N1842), .CI(N701));
ADDFXL inst_cellmath__203_0_I931 (.CO(N1880), .S(N1879), .A(N673), .B(N1875), .CI(N645));
ADDFX1 inst_cellmath__203_0_I932 (.CO(N1882), .S(N1881), .A(N729), .B(N1844), .CI(N757));
ADDFX1 inst_cellmath__203_0_I933 (.CO(N1884), .S(N1883), .A(N1848), .B(N1846), .CI(N1877));
ADDFX1 inst_cellmath__203_0_I934 (.CO(N1886), .S(N1885), .A(N1850), .B(N1879), .CI(N1881));
ADDFXL inst_cellmath__203_0_I935 (.CO(N1888), .S(N1887), .A(N1883), .B(N1852), .CI(N1854));
ADDFXL inst_cellmath__203_0_I936 (.CO(inst_cellmath__203_0_out1[26]), .S(inst_cellmath__203_0_out0[25]), .A(N1856), .B(N1885), .CI(N1887));
ADDHX1 inst_cellmath__203_0_I937 (.CO(N1892), .S(N1891), .A(N1860), .B(N1098));
ADDFX1 inst_cellmath__203_0_I938 (.CO(N1894), .S(N1893), .A(N1158), .B(N1128), .CI(N1891));
ADDFX1 inst_cellmath__203_0_I939 (.CO(N1896), .S(N1895), .A(N1248), .B(N1308), .CI(N1218));
ADDFX1 inst_cellmath__203_0_I940 (.CO(N1898), .S(N1897), .A(N1278), .B(N1188), .CI(N1864));
ADDFX1 inst_cellmath__203_0_I941 (.CO(N1900), .S(N1899), .A(N1868), .B(N1866), .CI(N1893));
ADDFX1 inst_cellmath__203_0_I942 (.CO(N1902), .S(N1901), .A(N1870), .B(N1895), .CI(N1897));
ADDFX1 inst_cellmath__203_0_I943 (.CO(N1904), .S(N1903), .A(N1899), .B(N1872), .CI(N1901));
ADDFX1 inst_cellmath__203_0_I944 (.CO(N1906), .S(N1905), .A(N5698), .B(N1874), .CI(N1876));
ADDFX1 inst_cellmath__203_0_I945 (.CO(N1908), .S(N1907), .A(N801), .B(N1903), .CI(N702));
ADDFX1 inst_cellmath__203_0_I946 (.CO(N1910), .S(N1909), .A(N730), .B(N674), .CI(N758));
ADDFXL inst_cellmath__203_0_I947 (.CO(N1912), .S(N1911), .A(N1878), .B(N1905), .CI(N1880));
ADDFX1 inst_cellmath__203_0_I948 (.CO(N1914), .S(N1913), .A(N1882), .B(N1907), .CI(N1909));
ADDFXL inst_cellmath__203_0_I949 (.CO(N1916), .S(N1915), .A(N1911), .B(N1884), .CI(N1886));
ADDFXL inst_cellmath__203_0_I950 (.CO(inst_cellmath__203_0_out1[27]), .S(inst_cellmath__203_0_out0[26]), .A(N1888), .B(N1913), .CI(N1915));
XNOR2X1 hap1_A_I1801 (.Y(N1919), .A(N1099), .B(N1249));
OR2XL hap1_A_I1802 (.Y(N1920), .A(N1099), .B(N1249));
ADDFX1 inst_cellmath__203_0_I952 (.CO(N1924), .S(N1923), .A(N1159), .B(N1129), .CI(N1189));
ADDFX1 inst_cellmath__203_0_I953 (.CO(N1926), .S(N1925), .A(N1279), .B(N1892), .CI(N1219));
ADDFX1 inst_cellmath__203_0_I954 (.CO(N1928), .S(N1927), .A(N1919), .B(N1309), .CI(N1894));
ADDFX1 inst_cellmath__203_0_I955 (.CO(N1930), .S(N1929), .A(N1923), .B(N1896), .CI(N1925));
ADDFX1 inst_cellmath__203_0_I956 (.CO(N1932), .S(N1931), .A(N1900), .B(N1898), .CI(N1927));
ADDFX1 inst_cellmath__203_0_I957 (.CO(N1934), .S(N1933), .A(N1902), .B(N1929), .CI(N1931));
ADDFX1 inst_cellmath__203_0_I958 (.CO(N1936), .S(N1935), .A(N803), .B(N1904), .CI(N703));
ADDFX1 inst_cellmath__203_0_I959 (.CO(N1938), .S(N1937), .A(N675), .B(N1933), .CI(N731));
ADDFX1 inst_cellmath__203_0_I960 (.CO(N1940), .S(N1939), .A(N759), .B(N1906), .CI(N1908));
ADDFX1 inst_cellmath__203_0_I961 (.CO(N1942), .S(N1941), .A(N1910), .B(N1935), .CI(N1937));
ADDFXL inst_cellmath__203_0_I962 (.CO(N1944), .S(N1943), .A(N1939), .B(N1912), .CI(N1914));
ADDFXL inst_cellmath__203_0_I963 (.CO(inst_cellmath__203_0_out1[28]), .S(inst_cellmath__203_0_out0[27]), .A(N1916), .B(N1941), .CI(N1943));
INVXL fap1_A_I1803 (.Y(N5435), .A(N5806));
ADDFX1 fap1_A_I1804 (.CO(N1948), .S(N1947), .A(N1160), .B(N1130), .CI(N5435));
ADDFX1 inst_cellmath__203_0_I965 (.CO(N1952), .S(N1951), .A(N1280), .B(N1190), .CI(N1250));
ADDFX1 inst_cellmath__203_0_I966 (.CO(N1954), .S(N1953), .A(N1310), .B(N1220), .CI(N1920));
ADDFX1 inst_cellmath__203_0_I967 (.CO(N1956), .S(N1955), .A(N1926), .B(N1924), .CI(N1951));
ADDFX1 inst_cellmath__203_0_I968 (.CO(N1958), .S(N1957), .A(N1953), .B(N1947), .CI(N1928));
ADDFX1 inst_cellmath__203_0_I969 (.CO(N1960), .S(N1959), .A(N1955), .B(N1930), .CI(N1957));
ADDFX1 inst_cellmath__203_0_I970 (.CO(N1962), .S(N1961), .A(N1959), .B(N1932), .CI(N5713));
ADDFX1 inst_cellmath__203_0_I971 (.CO(N1964), .S(N1963), .A(N805), .B(N1934), .CI(N704));
ADDFX1 inst_cellmath__203_0_I972 (.CO(N1966), .S(N1965), .A(N760), .B(N732), .CI(N1961));
ADDFX1 inst_cellmath__203_0_I973 (.CO(N1968), .S(N1967), .A(N1938), .B(N1936), .CI(N1963));
ADDFXL inst_cellmath__203_0_I974 (.CO(N1970), .S(N1969), .A(N1965), .B(N1940), .CI(N1942));
ADDFXL inst_cellmath__203_0_I975 (.CO(inst_cellmath__203_0_out1[29]), .S(inst_cellmath__203_0_out0[28]), .A(N1944), .B(N1967), .CI(N1969));
ADDFX1 inst_cellmath__203_0_I976 (.CO(N1974), .S(N1973), .A(N1131), .B(N5806), .CI(N1281));
ADDFX1 inst_cellmath__203_0_I977 (.CO(N1976), .S(N1975), .A(N1191), .B(N1161), .CI(N1221));
ADDFX1 inst_cellmath__203_0_I978 (.CO(N1978), .S(N1977), .A(N1251), .B(N1311), .CI(N1948));
ADDFX1 inst_cellmath__203_0_I979 (.CO(N1980), .S(N1979), .A(N1973), .B(N1952), .CI(N1954));
ADDFX1 inst_cellmath__203_0_I980 (.CO(N1982), .S(N1981), .A(N1977), .B(N1975), .CI(N1956));
ADDFX1 inst_cellmath__203_0_I981 (.CO(N1984), .S(N1983), .A(N1958), .B(N1979), .CI(N1981));
ADDFX1 inst_cellmath__203_0_I982 (.CO(N1986), .S(N1985), .A(N807), .B(N1960), .CI(N705));
ADDFX1 inst_cellmath__203_0_I983 (.CO(N1988), .S(N1987), .A(N1962), .B(N1983), .CI(N733));
ADDFX1 inst_cellmath__203_0_I984 (.CO(N1990), .S(N1989), .A(N1964), .B(N761), .CI(N1985));
ADDFX1 inst_cellmath__203_0_I985 (.CO(N1992), .S(N1991), .A(N1966), .B(N1987), .CI(N1968));
ADDFX1 inst_cellmath__203_0_I986 (.CO(inst_cellmath__203_0_out1[30]), .S(inst_cellmath__203_0_out0[29]), .A(N1970), .B(N1989), .CI(N1991));
INVXL fap1_A_I1805 (.Y(N5444), .A(N5842));
ADDFX1 fap1_A_I1806 (.CO(N1996), .S(N1995), .A(N1192), .B(N1162), .CI(N5444));
ADDFX1 inst_cellmath__203_0_I988 (.CO(N2000), .S(N1999), .A(N1312), .B(N1222), .CI(N1282));
ADDFX1 inst_cellmath__203_0_I989 (.CO(N2002), .S(N2001), .A(N1974), .B(N1252), .CI(N1976));
ADDFX1 inst_cellmath__203_0_I990 (.CO(N2004), .S(N2003), .A(N1995), .B(N1999), .CI(N1978));
ADDFX1 inst_cellmath__203_0_I991 (.CO(N2006), .S(N2005), .A(N2001), .B(N1980), .CI(N2003));
ADDFX1 inst_cellmath__203_0_I992 (.CO(N2008), .S(N2007), .A(N2005), .B(N1982), .CI(N5731));
ADDFX1 inst_cellmath__203_0_I993 (.CO(N2010), .S(N2009), .A(N809), .B(N1984), .CI(N734));
ADDFX1 inst_cellmath__203_0_I994 (.CO(N2012), .S(N2011), .A(N762), .B(N2007), .CI(N1986));
ADDFX1 inst_cellmath__203_0_I995 (.CO(N2014), .S(N2013), .A(N2009), .B(N1988), .CI(N1990));
ADDFX1 inst_cellmath__203_0_I996 (.CO(inst_cellmath__203_0_out1[31]), .S(inst_cellmath__203_0_out0[30]), .A(N1992), .B(N2011), .CI(N2013));
ADDFX1 inst_cellmath__203_0_I997 (.CO(N2018), .S(N2017), .A(N1163), .B(N5842), .CI(N1313));
ADDFX1 inst_cellmath__203_0_I998 (.CO(N2020), .S(N2019), .A(N1223), .B(N1193), .CI(N1253));
ADDFX1 inst_cellmath__203_0_I999 (.CO(N2022), .S(N2021), .A(N1996), .B(N1283), .CI(N2000));
ADDFX1 inst_cellmath__203_0_I1000 (.CO(N2024), .S(N2023), .A(N2019), .B(N2017), .CI(N2002));
ADDFX1 inst_cellmath__203_0_I1001 (.CO(N2026), .S(N2025), .A(N2004), .B(N2021), .CI(N2023));
ADDFX1 inst_cellmath__203_0_I1002 (.CO(N2028), .S(N2027), .A(N2025), .B(N2006), .CI(N811));
ADDFX1 inst_cellmath__203_0_I1003 (.CO(N2030), .S(N2029), .A(N735), .B(N2008), .CI(N763));
ADDFX1 inst_cellmath__203_0_I1004 (.CO(N2032), .S(N2031), .A(N2027), .B(N2010), .CI(N2012));
ADDFX1 inst_cellmath__203_0_I1005 (.CO(inst_cellmath__203_0_out1[32]), .S(inst_cellmath__203_0_out0[31]), .A(N2014), .B(N2029), .CI(N2031));
INVXL fap1_A_I1807 (.Y(N5453), .A(N5868));
ADDFX1 fap1_A_I1808 (.CO(N2036), .S(N2035), .A(N1224), .B(N1194), .CI(N5453));
ADDFX1 inst_cellmath__203_0_I1007 (.CO(N2040), .S(N2039), .A(N1314), .B(N1254), .CI(N1284));
ADDFX1 inst_cellmath__203_0_I1008 (.CO(N2042), .S(N2041), .A(N2020), .B(N2018), .CI(N2035));
ADDFX1 inst_cellmath__203_0_I1009 (.CO(N2044), .S(N2043), .A(N2022), .B(N2039), .CI(N2024));
ADDFX1 inst_cellmath__203_0_I1010 (.CO(N2046), .S(N2045), .A(N2026), .B(N2041), .CI(N2043));
ADDFX1 inst_cellmath__203_0_I1011 (.CO(N2048), .S(N2047), .A(N813), .B(N5747), .CI(N2045));
ADDFX1 inst_cellmath__203_0_I1012 (.CO(N2050), .S(N2049), .A(N2028), .B(N764), .CI(N2047));
ADDFXL inst_cellmath__203_0_I1013 (.CO(inst_cellmath__203_0_out0[33]), .S(inst_cellmath__203_0_out0[32]), .A(N2049), .B(N2030), .CI(N2032));
ADDFX1 inst_cellmath__203_0_I1014 (.CO(N2054), .S(N2053), .A(N1195), .B(N5868), .CI(N1225));
ADDFX1 inst_cellmath__203_0_I1015 (.CO(N2056), .S(N2055), .A(N1285), .B(N1255), .CI(N1315));
ADDFX1 inst_cellmath__203_0_I1016 (.CO(N2058), .S(N2057), .A(N2040), .B(N2036), .CI(N2053));
ADDFX1 inst_cellmath__203_0_I1017 (.CO(N2060), .S(N2059), .A(N2042), .B(N2055), .CI(N2057));
ADDFX1 inst_cellmath__203_0_I1018 (.CO(N2062), .S(N2061), .A(N2059), .B(N2044), .CI(N2046));
ADDFX1 inst_cellmath__203_0_I1019 (.CO(N2064), .S(N2063), .A(N765), .B(N815), .CI(N2061));
ADDFX1 inst_cellmath__203_0_I1020 (.CO(inst_cellmath__203_0_out0[34]), .S(inst_cellmath__203_0_out1[33]), .A(N2063), .B(N2048), .CI(N2050));
INVXL fap1_A_I1809 (.Y(N5462), .A(N5896));
ADDFX1 fap1_A_I1810 (.CO(N2068), .S(N2067), .A(N1256), .B(N1226), .CI(N5462));
ADDFX1 inst_cellmath__203_0_I1022 (.CO(N2072), .S(N2071), .A(N1316), .B(N1286), .CI(N2054));
ADDFX1 inst_cellmath__203_0_I1023 (.CO(N2074), .S(N2073), .A(N2067), .B(N2056), .CI(N2058));
ADDFX1 inst_cellmath__203_0_I1024 (.CO(N2076), .S(N2075), .A(N2060), .B(N2071), .CI(N2073));
ADDFX1 inst_cellmath__203_0_I1025 (.CO(N2078), .S(N2077), .A(N817), .B(N2075), .CI(N5763));
ADDFX1 inst_cellmath__203_0_I1026 (.CO(inst_cellmath__203_0_out0[35]), .S(inst_cellmath__203_0_out1[34]), .A(N2077), .B(N2062), .CI(N2064));
ADDFX1 inst_cellmath__203_0_I1027 (.CO(N2082), .S(N2081), .A(N1227), .B(N5896), .CI(N1257));
ADDFX1 inst_cellmath__203_0_I1028 (.CO(N2084), .S(N2083), .A(N1317), .B(N1287), .CI(N2068));
ADDFX1 inst_cellmath__203_0_I1029 (.CO(N2086), .S(N2085), .A(N2072), .B(N2081), .CI(N2083));
ADDFX1 inst_cellmath__203_0_I1030 (.CO(N2088), .S(N2087), .A(N2085), .B(N2074), .CI(N2076));
ADDFX1 inst_cellmath__203_0_I1031 (.CO(inst_cellmath__203_0_out0[36]), .S(inst_cellmath__203_0_out1[35]), .A(N2087), .B(N819), .CI(N2078));
INVXL fap1_A_I1811 (.Y(N5471), .A(N5924));
ADDFX1 fap1_A_I1812 (.CO(N2092), .S(N2091), .A(N1288), .B(N1258), .CI(N5471));
ADDFX1 inst_cellmath__203_0_I1033 (.CO(N2096), .S(N2095), .A(N2082), .B(N1318), .CI(N2091));
ADDFX1 inst_cellmath__203_0_I1034 (.CO(N2098), .S(N2097), .A(N2095), .B(N2084), .CI(N2086));
ADDFX1 inst_cellmath__203_0_I1035 (.CO(inst_cellmath__203_0_out0[37]), .S(inst_cellmath__203_0_out1[36]), .A(N1366), .B(N2097), .CI(N2088));
ADDFX1 inst_cellmath__203_0_I1036 (.CO(N2102), .S(N2101), .A(N1259), .B(N5924), .CI(N1289));
ADDFX1 inst_cellmath__203_0_I1037 (.CO(N2104), .S(N2103), .A(N2092), .B(N1319), .CI(N2101));
ADDFX1 inst_cellmath__203_0_I1038 (.CO(inst_cellmath__203_0_out0[38]), .S(inst_cellmath__203_0_out1[37]), .A(N2103), .B(N2096), .CI(N2098));
ADDFX1 inst_cellmath__203_0_I1039 (.CO(N2108), .S(N2107), .A(N1290), .B(N5947), .CI(N1320));
ADDFX1 inst_cellmath__203_0_I1040 (.CO(inst_cellmath__203_0_out0[39]), .S(inst_cellmath__203_0_out1[38]), .A(N2107), .B(N2102), .CI(N2104));
INVXL inst_cellmath__203_0_I1041 (.Y(N2111), .A(N2112));
ADDFX1 inst_cellmath__203_0_I1042 (.CO(inst_cellmath__203_0_out0[40]), .S(inst_cellmath__203_0_out1[39]), .A(N1321), .B(N2111), .CI(N2108));
ADDFX1 inst_cellmath__203_0_I1043 (.CO(inst_cellmath__203_0_out0[41]), .S(inst_cellmath__203_0_out1[40]), .A(N2112), .B(N5970), .CI(N1322));
INVXL inst_cellmath__203_0_I1044 (.Y(inst_cellmath__203_0_out1[41]), .A(inst_cellmath__203_0_out0[42]));
assign inst_cellmath__203_0_out0[0] = 1'B0;
assign inst_cellmath__203_0_out0[43] = 1'B0;
assign inst_cellmath__203_0_out0[44] = 1'B0;
assign inst_cellmath__203_0_out0[45] = 1'B0;
assign inst_cellmath__203_0_out0[46] = 1'B0;
assign inst_cellmath__203_0_out1[43] = 1'B1;
assign inst_cellmath__203_0_out1[44] = 1'B1;
assign inst_cellmath__203_0_out1[45] = 1'B1;
assign inst_cellmath__203_0_out1[46] = 1'B1;
endmodule

module cynw_cm_float_sin_inst_cellmath__201_0_bdw1946085813_bdw (
	inst_cellmath__201_0_out0,
	inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1,
	inst_cellmath__201_0_in2
	); /* architecture "gate_level" */ 
output [49:0] inst_cellmath__201_0_out0;
input [46:0] inst_cellmath__201_0_in0,
	inst_cellmath__201_0_in1;
input [72:43] inst_cellmath__201_0_in2;
wire [46:0] inst_cellmath__203__W1;
wire N989,N991,N992,N993,N994,N995,N996 
	,N997,N998,N999,N1000,N1001,N1002,N1003,N1004 
	,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012 
	,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020 
	,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028 
	,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036 
	,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044 
	,N1045,N1046,N1047,N1048,N1049,N1053,N1054,N1055 
	,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063 
	,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071 
	,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079 
	,N1080,N1081,N1082,N1083,N1084,N1085,N1088,N1092 
	,N1093,N1100,N1110,N1114,N1115,N1128,N1144,N1164 
	,N1168,N1192,N1194,N1220,N1254,N1256,N1260,N1261 
	,N1292,N1326,N1350,N1353,N1356,N1359,N1362,N1365 
	,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389 
	,N1392,N1395,N1413,N1415,N1416,N1417,N1418,N1419 
	,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427 
	,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435 
	,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443 
	,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451 
	,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459 
	,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467 
	,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475 
	,N1476,N1480,N1484,N1485,N1488,N1489,N1492,N1493 
	,N1496,N1497,N1500,N1501,N1504,N1505,N1508,N1509 
	,N1512,N1513,N1516,N1517,N1520,N1521,N1532,N1533 
	,N1536,N1537,N1548,N1549,N1552,N1553,N1564,N1565 
	,N1572,N1607,N1609,N1610,N1611,N1612,N1613,N1614 
	,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622 
	,N1623,N1624,N1625,N1626,N1627,N1628,N1633,N1635 
	,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644 
	,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652 
	,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676 
	,N1693,N1695,N1697,N1699,N1739,N1742,N1745,N1748 
	,N1751,N1754,N1757,N1760,N1763,N1766,N1769,N1772 
	,N1775,N1778,N1781,N1784,N1787,N1790,N1793,N1802 
	,N1805,N1814,N1817,N1826,N1829,N1848,N1849,N1851 
	,N1852,N1854,N1855,N1857,N1858,N1860,N1861,N1863 
	,N1864,N1866,N1867,N1869,N1870,N1872,N1873,N1875 
	,N1876,N1878,N1879,N1881,N1882,N1884,N1885,N1887 
	,N1888,N1890,N1891,N1893,N1894,N1896,N1897,N1899 
	,N1900,N1902,N1903,N1907,N2056,N2058,N2067,N2069 
	,N2085,N2087,N2096,N2098,N2114,N2116,N2125,N2127 
	,N2143,N2308,N2309,N2322,N2323,N2333,N2334,N2352 
	,N2353,N2369,N2386,N2389,N2398,N2420,N2428,N2436 
	,N2443,N2452,N2454,N2455,N2460,N2462,N2463,N2468 
	,N2470,N2471,N2477,N2478,N2479,N2480,N2483,N2484 
	,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492 
	,N2493,N2494,N2496,N2524,N2531,N2538,N2545,N2552 
	,N2559,N3749;
INVXL inst_cellmath__201_0_I102 (.Y(inst_cellmath__203__W1[46]), .A(inst_cellmath__201_0_in0[46]));
INVXL inst_cellmath__201_0_I243 (.Y(N989), .A(inst_cellmath__201_0_in1[46]));
ADDHX1 inst_cellmath__201_0_I245 (.CO(N992), .S(N991), .A(inst_cellmath__201_0_in2[43]), .B(inst_cellmath__201_0_in1[18]));
ADDFX1 inst_cellmath__201_0_I246 (.CO(N994), .S(N993), .A(inst_cellmath__201_0_in1[19]), .B(inst_cellmath__201_0_in2[44]), .CI(inst_cellmath__201_0_in0[19]));
ADDFX1 inst_cellmath__201_0_I247 (.CO(N996), .S(N995), .A(inst_cellmath__201_0_in1[20]), .B(inst_cellmath__201_0_in2[45]), .CI(inst_cellmath__201_0_in0[20]));
ADDFX1 inst_cellmath__201_0_I248 (.CO(N998), .S(N997), .A(inst_cellmath__201_0_in1[21]), .B(inst_cellmath__201_0_in2[46]), .CI(inst_cellmath__201_0_in0[21]));
ADDFX1 inst_cellmath__201_0_I249 (.CO(N1000), .S(N999), .A(inst_cellmath__201_0_in1[22]), .B(inst_cellmath__201_0_in2[47]), .CI(inst_cellmath__201_0_in0[22]));
ADDFHXL inst_cellmath__201_0_I250 (.CO(N1002), .S(N1001), .A(inst_cellmath__201_0_in1[23]), .B(inst_cellmath__201_0_in2[48]), .CI(inst_cellmath__201_0_in0[23]));
ADDFX1 inst_cellmath__201_0_I251 (.CO(N1004), .S(N1003), .A(inst_cellmath__201_0_in1[24]), .B(inst_cellmath__201_0_in2[49]), .CI(inst_cellmath__201_0_in0[24]));
ADDFX1 inst_cellmath__201_0_I252 (.CO(N1006), .S(N1005), .A(inst_cellmath__201_0_in1[25]), .B(inst_cellmath__201_0_in2[50]), .CI(inst_cellmath__201_0_in0[25]));
ADDFXL inst_cellmath__201_0_I253 (.CO(N1008), .S(N1007), .A(inst_cellmath__201_0_in1[26]), .B(inst_cellmath__201_0_in2[51]), .CI(inst_cellmath__201_0_in0[26]));
ADDFX1 inst_cellmath__201_0_I254 (.CO(N1010), .S(N1009), .A(inst_cellmath__201_0_in1[27]), .B(inst_cellmath__201_0_in2[52]), .CI(inst_cellmath__201_0_in0[27]));
ADDFX1 inst_cellmath__201_0_I255 (.CO(N1012), .S(N1011), .A(inst_cellmath__201_0_in1[28]), .B(inst_cellmath__201_0_in2[53]), .CI(inst_cellmath__201_0_in0[28]));
ADDFX1 inst_cellmath__201_0_I256 (.CO(N1014), .S(N1013), .A(inst_cellmath__201_0_in1[29]), .B(inst_cellmath__201_0_in2[54]), .CI(inst_cellmath__201_0_in0[29]));
ADDFX1 inst_cellmath__201_0_I257 (.CO(N1016), .S(N1015), .A(inst_cellmath__201_0_in1[30]), .B(inst_cellmath__201_0_in2[55]), .CI(inst_cellmath__201_0_in0[30]));
ADDFX1 inst_cellmath__201_0_I258 (.CO(N1018), .S(N1017), .A(inst_cellmath__201_0_in1[31]), .B(inst_cellmath__201_0_in2[56]), .CI(inst_cellmath__201_0_in0[31]));
ADDFX1 inst_cellmath__201_0_I259 (.CO(N1020), .S(N1019), .A(inst_cellmath__201_0_in0[32]), .B(inst_cellmath__201_0_in2[57]), .CI(inst_cellmath__201_0_in1[32]));
ADDFX1 inst_cellmath__201_0_I260 (.CO(N1022), .S(N1021), .A(inst_cellmath__201_0_in0[33]), .B(inst_cellmath__201_0_in2[58]), .CI(inst_cellmath__201_0_in1[33]));
ADDFX1 inst_cellmath__201_0_I261 (.CO(N1024), .S(N1023), .A(inst_cellmath__201_0_in1[34]), .B(inst_cellmath__201_0_in2[59]), .CI(inst_cellmath__201_0_in0[34]));
ADDFX1 inst_cellmath__201_0_I262 (.CO(N1026), .S(N1025), .A(inst_cellmath__201_0_in0[35]), .B(inst_cellmath__201_0_in2[60]), .CI(inst_cellmath__201_0_in1[35]));
ADDFX1 inst_cellmath__201_0_I263 (.CO(N1028), .S(N1027), .A(inst_cellmath__201_0_in1[36]), .B(inst_cellmath__201_0_in2[61]), .CI(inst_cellmath__201_0_in0[36]));
ADDFX1 inst_cellmath__201_0_I264 (.CO(N1030), .S(N1029), .A(inst_cellmath__201_0_in1[37]), .B(inst_cellmath__201_0_in2[62]), .CI(inst_cellmath__201_0_in0[37]));
ADDFX1 inst_cellmath__201_0_I265 (.CO(N1032), .S(N1031), .A(inst_cellmath__201_0_in1[38]), .B(inst_cellmath__201_0_in2[63]), .CI(inst_cellmath__201_0_in0[38]));
ADDFX1 inst_cellmath__201_0_I266 (.CO(N1034), .S(N1033), .A(inst_cellmath__201_0_in1[39]), .B(inst_cellmath__201_0_in2[64]), .CI(inst_cellmath__201_0_in0[39]));
ADDFX1 inst_cellmath__201_0_I267 (.CO(N1036), .S(N1035), .A(inst_cellmath__201_0_in1[40]), .B(inst_cellmath__201_0_in2[65]), .CI(inst_cellmath__201_0_in0[40]));
ADDFX1 inst_cellmath__201_0_I268 (.CO(N1038), .S(N1037), .A(inst_cellmath__201_0_in1[41]), .B(inst_cellmath__201_0_in2[66]), .CI(inst_cellmath__201_0_in0[41]));
ADDFX1 inst_cellmath__201_0_I269 (.CO(N1040), .S(N1039), .A(inst_cellmath__201_0_in0[42]), .B(inst_cellmath__201_0_in1[42]), .CI(inst_cellmath__201_0_in2[67]));
ADDFX1 inst_cellmath__201_0_I270 (.CO(N1042), .S(N1041), .A(inst_cellmath__201_0_in0[43]), .B(inst_cellmath__201_0_in1[43]), .CI(inst_cellmath__201_0_in2[68]));
ADDFX1 inst_cellmath__201_0_I271 (.CO(N1044), .S(N1043), .A(inst_cellmath__201_0_in0[44]), .B(inst_cellmath__201_0_in1[44]), .CI(inst_cellmath__201_0_in2[69]));
ADDFX1 inst_cellmath__201_0_I272 (.CO(N1046), .S(N1045), .A(inst_cellmath__201_0_in0[45]), .B(inst_cellmath__201_0_in1[45]), .CI(inst_cellmath__201_0_in2[70]));
ADDFX1 inst_cellmath__201_0_I273 (.CO(N1048), .S(N1047), .A(inst_cellmath__203__W1[46]), .B(N989), .CI(inst_cellmath__201_0_in2[71]));
INVXL inst_cellmath__201_0_I274 (.Y(N1049), .A(inst_cellmath__201_0_in2[72]));
NAND2XL inst_cellmath__201_0_I275 (.Y(N1053), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
NOR2XL inst_cellmath__201_0_I276 (.Y(N1054), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NAND2XL inst_cellmath__201_0_I277 (.Y(N1055), .A(inst_cellmath__201_0_in1[1]), .B(inst_cellmath__201_0_in0[1]));
NOR2XL inst_cellmath__201_0_I278 (.Y(N1056), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NAND2XL inst_cellmath__201_0_I279 (.Y(N1057), .A(inst_cellmath__201_0_in1[2]), .B(inst_cellmath__201_0_in0[2]));
NOR2XL inst_cellmath__201_0_I280 (.Y(N1058), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NAND2XL inst_cellmath__201_0_I281 (.Y(N1059), .A(inst_cellmath__201_0_in1[3]), .B(inst_cellmath__201_0_in0[3]));
NOR2XL inst_cellmath__201_0_I282 (.Y(N1060), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NAND2XL inst_cellmath__201_0_I283 (.Y(N1061), .A(inst_cellmath__201_0_in1[4]), .B(inst_cellmath__201_0_in0[4]));
NOR2XL inst_cellmath__201_0_I284 (.Y(N1062), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NAND2XL inst_cellmath__201_0_I285 (.Y(N1063), .A(inst_cellmath__201_0_in1[5]), .B(inst_cellmath__201_0_in0[5]));
NOR2XL inst_cellmath__201_0_I286 (.Y(N1064), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NAND2XL inst_cellmath__201_0_I287 (.Y(N1065), .A(inst_cellmath__201_0_in1[6]), .B(inst_cellmath__201_0_in0[6]));
NOR2XL inst_cellmath__201_0_I288 (.Y(N1066), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NAND2XL inst_cellmath__201_0_I289 (.Y(N1067), .A(inst_cellmath__201_0_in1[7]), .B(inst_cellmath__201_0_in0[7]));
NOR2XL inst_cellmath__201_0_I290 (.Y(N1068), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NAND2XL inst_cellmath__201_0_I291 (.Y(N1069), .A(inst_cellmath__201_0_in1[8]), .B(inst_cellmath__201_0_in0[8]));
NOR2XL inst_cellmath__201_0_I292 (.Y(N1070), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NAND2XL inst_cellmath__201_0_I293 (.Y(N1071), .A(inst_cellmath__201_0_in1[9]), .B(inst_cellmath__201_0_in0[9]));
NOR2XL inst_cellmath__201_0_I294 (.Y(N1072), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NAND2X1 inst_cellmath__201_0_I295 (.Y(N1073), .A(inst_cellmath__201_0_in1[10]), .B(inst_cellmath__201_0_in0[10]));
NOR2XL inst_cellmath__201_0_I296 (.Y(N1074), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NAND2XL inst_cellmath__201_0_I297 (.Y(N1075), .A(inst_cellmath__201_0_in1[11]), .B(inst_cellmath__201_0_in0[11]));
NOR2XL inst_cellmath__201_0_I298 (.Y(N1076), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NAND2XL inst_cellmath__201_0_I299 (.Y(N1077), .A(inst_cellmath__201_0_in1[12]), .B(inst_cellmath__201_0_in0[12]));
NOR2XL inst_cellmath__201_0_I300 (.Y(N1078), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NAND2X1 inst_cellmath__201_0_I301 (.Y(N1079), .A(inst_cellmath__201_0_in1[13]), .B(inst_cellmath__201_0_in0[13]));
NOR2XL inst_cellmath__201_0_I302 (.Y(N1080), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NAND2XL inst_cellmath__201_0_I303 (.Y(N1081), .A(inst_cellmath__201_0_in1[14]), .B(inst_cellmath__201_0_in0[14]));
NOR2XL inst_cellmath__201_0_I304 (.Y(N1082), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NAND2XL inst_cellmath__201_0_I305 (.Y(N1083), .A(inst_cellmath__201_0_in1[15]), .B(inst_cellmath__201_0_in0[15]));
NOR2XL inst_cellmath__201_0_I306 (.Y(N1084), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
NAND2XL inst_cellmath__201_0_I307 (.Y(N1085), .A(inst_cellmath__201_0_in1[16]), .B(inst_cellmath__201_0_in0[16]));
AOI21XL inst_cellmath__201_0_I310 (.Y(N1088), .A0(N1055), .A1(N1053), .B0(N1054));
AOI21XL inst_cellmath__201_0_I314 (.Y(N1092), .A0(N1059), .A1(N1056), .B0(N1058));
NAND2XL inst_cellmath__201_0_I315 (.Y(N1093), .A(N1059), .B(N1057));
OAI21XL inst_cellmath__201_0_I322 (.Y(N1100), .A0(N1093), .A1(N1088), .B0(N1092));
AOI21XL inst_cellmath__201_0_I332 (.Y(N1110), .A0(N1061), .A1(N1100), .B0(N1060));
AOI21XL inst_cellmath__201_0_I336 (.Y(N1114), .A0(N1065), .A1(N1062), .B0(N1064));
NAND2XL inst_cellmath__201_0_I337 (.Y(N1115), .A(N1065), .B(N1063));
OAI21XL inst_cellmath__201_0_I350 (.Y(N1128), .A0(N1115), .A1(N1110), .B0(N1114));
AOI21XL inst_cellmath__201_0_I366 (.Y(N1144), .A0(N1067), .A1(N1128), .B0(N1066));
INVXL inst_cellmath__201_0_I1260 (.Y(N2308), .A(N1068));
INVXL inst_cellmath__201_0_I1261 (.Y(N2309), .A(N1069));
OAI21X1 inst_cellmath__201_0_I386 (.Y(N1164), .A0(N2309), .A1(N1144), .B0(N2308));
AOI21XL inst_cellmath__201_0_I390 (.Y(N1168), .A0(N1073), .A1(N1070), .B0(N1072));
INVXL inst_cellmath__201_0_I1274 (.Y(N2322), .A(N1168));
AND2XL inst_cellmath__201_0_I1463 (.Y(N2323), .A(N1073), .B(N1071));
AOI21XL inst_cellmath__201_0_I414 (.Y(N1192), .A0(N1071), .A1(N1164), .B0(N1070));
AOI21X2 inst_cellmath__201_0_I416 (.Y(N1194), .A0(N2323), .A1(N1164), .B0(N2322));
INVXL inst_cellmath__201_0_I1285 (.Y(N2333), .A(N1074));
INVXL inst_cellmath__201_0_I1286 (.Y(N2334), .A(N1075));
OAI21X2 inst_cellmath__201_0_I442 (.Y(N1220), .A0(N2334), .A1(N1194), .B0(N2333));
AO21XL inst_cellmath__201_0_I1465 (.Y(N2352), .A0(N1079), .A1(N1076), .B0(N1078));
AND2X1 inst_cellmath__201_0_I1451 (.Y(N2353), .A(N1077), .B(N1079));
AOI21XL inst_cellmath__201_0_I476 (.Y(N1254), .A0(N1077), .A1(N1220), .B0(N1076));
AOI21X4 inst_cellmath__201_0_I478 (.Y(N1256), .A0(N2353), .A1(N1220), .B0(N2352));
INVXL inst_cellmath__201_0_I1321 (.Y(N2369), .A(N1081));
AOI21XL inst_cellmath__201_0_I482 (.Y(N1260), .A0(N1083), .A1(N1080), .B0(N1082));
NAND2XL inst_cellmath__201_0_I483 (.Y(N1261), .A(N1083), .B(N1081));
OAI21X2 inst_cellmath__201_0_I514 (.Y(N1292), .A0(N1261), .A1(N1256), .B0(N1260));
NOR2BX1 andori2bb1_A_I2447 (.Y(N2524), .AN(N1057), .B(N1088));
NOR2XL andori2bb1_A_I1569 (.Y(N2386), .A(N2524), .B(N1056));
NOR2BX1 andori2bb1_A_I2448 (.Y(N2531), .AN(N1063), .B(N1110));
NOR2XL andori2bb1_A_I1571 (.Y(N2389), .A(N2531), .B(N1062));
NOR2XL andori2bb1_A_I1572 (.Y(N2538), .A(N2369), .B(N1256));
NOR2XL andori2bb1_A_I1573 (.Y(N2398), .A(N2538), .B(N1080));
AOI21X2 inst_cellmath__201_0_I548 (.Y(N1326), .A0(N1085), .A1(N1292), .B0(N1084));
NAND2BXL inst_cellmath__201_0_I572 (.Y(N1350), .AN(N1054), .B(N1055));
NAND2BXL inst_cellmath__201_0_I575 (.Y(N1353), .AN(N1056), .B(N1057));
NAND2BXL inst_cellmath__201_0_I578 (.Y(N1356), .AN(N1058), .B(N1059));
NAND2BXL inst_cellmath__201_0_I581 (.Y(N1359), .AN(N1060), .B(N1061));
NAND2BXL inst_cellmath__201_0_I584 (.Y(N1362), .AN(N1062), .B(N1063));
NAND2BXL inst_cellmath__201_0_I587 (.Y(N1365), .AN(N1064), .B(N1065));
NAND2BXL inst_cellmath__201_0_I590 (.Y(N1368), .AN(N1066), .B(N1067));
NAND2BXL inst_cellmath__201_0_I593 (.Y(N1371), .AN(N1068), .B(N1069));
NAND2BXL inst_cellmath__201_0_I596 (.Y(N1374), .AN(N1070), .B(N1071));
NAND2BXL inst_cellmath__201_0_I599 (.Y(N1377), .AN(N1072), .B(N1073));
NAND2BXL inst_cellmath__201_0_I602 (.Y(N1380), .AN(N1074), .B(N1075));
NAND2BXL inst_cellmath__201_0_I605 (.Y(N1383), .AN(N1076), .B(N1077));
NAND2BXL inst_cellmath__201_0_I608 (.Y(N1386), .AN(N1078), .B(N1079));
NAND2BXL inst_cellmath__201_0_I611 (.Y(N1389), .AN(N1080), .B(N1081));
NAND2BXL inst_cellmath__201_0_I614 (.Y(N1392), .AN(N1082), .B(N1083));
NAND2BXL inst_cellmath__201_0_I617 (.Y(N1395), .AN(N1084), .B(N1085));
XOR2XL inst_cellmath__201_0_I618 (.Y(inst_cellmath__201_0_out0[0]), .A(inst_cellmath__201_0_in0[0]), .B(inst_cellmath__201_0_in1[0]));
XOR2XL inst_cellmath__201_0_I1471 (.Y(inst_cellmath__201_0_out0[1]), .A(N1053), .B(N1350));
XNOR2X1 inst_cellmath__201_0_I620 (.Y(inst_cellmath__201_0_out0[2]), .A(N1088), .B(N1353));
XNOR2X1 inst_cellmath__201_0_I621 (.Y(inst_cellmath__201_0_out0[3]), .A(N2386), .B(N1356));
XOR2XL inst_cellmath__201_0_I1472 (.Y(inst_cellmath__201_0_out0[4]), .A(N1100), .B(N1359));
XNOR2X1 inst_cellmath__201_0_I623 (.Y(inst_cellmath__201_0_out0[5]), .A(N1110), .B(N1362));
XNOR2X1 inst_cellmath__201_0_I624 (.Y(inst_cellmath__201_0_out0[6]), .A(N2389), .B(N1365));
XOR2XL inst_cellmath__201_0_I1473 (.Y(inst_cellmath__201_0_out0[7]), .A(N1128), .B(N1368));
XNOR2X1 inst_cellmath__201_0_I626 (.Y(inst_cellmath__201_0_out0[8]), .A(N1144), .B(N1371));
XOR2XL inst_cellmath__201_0_I1474 (.Y(inst_cellmath__201_0_out0[9]), .A(N1164), .B(N1374));
XNOR2X1 inst_cellmath__201_0_I628 (.Y(inst_cellmath__201_0_out0[10]), .A(N1192), .B(N1377));
XNOR2X1 inst_cellmath__201_0_I629 (.Y(inst_cellmath__201_0_out0[11]), .A(N1194), .B(N1380));
XOR2XL inst_cellmath__201_0_I1475 (.Y(inst_cellmath__201_0_out0[12]), .A(N1220), .B(N1383));
XNOR2X1 inst_cellmath__201_0_I631 (.Y(inst_cellmath__201_0_out0[13]), .A(N1254), .B(N1386));
XNOR2X1 inst_cellmath__201_0_I632 (.Y(inst_cellmath__201_0_out0[14]), .A(N1256), .B(N1389));
XNOR2X1 inst_cellmath__201_0_I633 (.Y(inst_cellmath__201_0_out0[15]), .A(N2398), .B(N1392));
XOR2XL inst_cellmath__201_0_I1476 (.Y(inst_cellmath__201_0_out0[16]), .A(N1292), .B(N1395));
INVX2 inst_cellmath__201_0_I635 (.Y(N1413), .A(N1326));
NOR2XL inst_cellmath__201_0_I636 (.Y(N1415), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NAND2XL inst_cellmath__201_0_I637 (.Y(N1416), .A(inst_cellmath__201_0_in1[17]), .B(inst_cellmath__201_0_in0[17]));
NOR2XL inst_cellmath__201_0_I638 (.Y(N1417), .A(N991), .B(inst_cellmath__201_0_in0[18]));
NAND2XL inst_cellmath__201_0_I639 (.Y(N1418), .A(N991), .B(inst_cellmath__201_0_in0[18]));
NOR2X1 inst_cellmath__201_0_I640 (.Y(N1419), .A(N992), .B(N993));
NAND2X2 inst_cellmath__201_0_I641 (.Y(N1420), .A(N992), .B(N993));
NOR2X2 inst_cellmath__201_0_I642 (.Y(N1421), .A(N994), .B(N995));
NAND2X2 inst_cellmath__201_0_I643 (.Y(N1422), .A(N994), .B(N995));
NOR2X1 inst_cellmath__201_0_I644 (.Y(N1423), .A(N996), .B(N997));
NAND2X4 inst_cellmath__201_0_I645 (.Y(N1424), .A(N996), .B(N997));
NOR2X2 inst_cellmath__201_0_I646 (.Y(N1425), .A(N998), .B(N999));
NAND2X2 inst_cellmath__201_0_I647 (.Y(N1426), .A(N998), .B(N999));
NOR2X1 inst_cellmath__201_0_I648 (.Y(N1427), .A(N1000), .B(N1001));
NAND2X4 inst_cellmath__201_0_I649 (.Y(N1428), .A(N1000), .B(N1001));
NOR2X4 inst_cellmath__201_0_I650 (.Y(N1429), .A(N1002), .B(N1003));
NAND2X2 inst_cellmath__201_0_I651 (.Y(N1430), .A(N1002), .B(N1003));
NOR2X1 inst_cellmath__201_0_I652 (.Y(N1431), .A(N1004), .B(N1005));
NAND2X4 inst_cellmath__201_0_I653 (.Y(N1432), .A(N1004), .B(N1005));
NOR2X1 inst_cellmath__201_0_I654 (.Y(N1433), .A(N1006), .B(N1007));
NAND2X1 inst_cellmath__201_0_I655 (.Y(N1434), .A(N1006), .B(N1007));
NOR2X1 inst_cellmath__201_0_I656 (.Y(N1435), .A(N1008), .B(N1009));
NAND2X4 inst_cellmath__201_0_I657 (.Y(N1436), .A(N1008), .B(N1009));
NOR2X1 inst_cellmath__201_0_I658 (.Y(N1437), .A(N1010), .B(N1011));
NAND2X1 inst_cellmath__201_0_I659 (.Y(N1438), .A(N1010), .B(N1011));
NOR2XL inst_cellmath__201_0_I660 (.Y(N1439), .A(N1012), .B(N1013));
NAND2X2 inst_cellmath__201_0_I661 (.Y(N1440), .A(N1012), .B(N1013));
NOR2XL inst_cellmath__201_0_I662 (.Y(N1441), .A(N1014), .B(N1015));
NAND2XL inst_cellmath__201_0_I663 (.Y(N1442), .A(N1014), .B(N1015));
NOR2XL inst_cellmath__201_0_I664 (.Y(N1443), .A(N1016), .B(N1017));
NAND2XL inst_cellmath__201_0_I665 (.Y(N1444), .A(N1016), .B(N1017));
NOR2XL inst_cellmath__201_0_I666 (.Y(N1445), .A(N1018), .B(N1019));
NAND2XL inst_cellmath__201_0_I667 (.Y(N1446), .A(N1018), .B(N1019));
NOR2XL inst_cellmath__201_0_I668 (.Y(N1447), .A(N1021), .B(N1020));
NAND2XL inst_cellmath__201_0_I669 (.Y(N1448), .A(N1021), .B(N1020));
NOR2XL inst_cellmath__201_0_I670 (.Y(N1449), .A(N1023), .B(N1022));
NAND2XL inst_cellmath__201_0_I671 (.Y(N1450), .A(N1023), .B(N1022));
NOR2XL inst_cellmath__201_0_I672 (.Y(N1451), .A(N1024), .B(N1025));
NAND2XL inst_cellmath__201_0_I673 (.Y(N1452), .A(N1024), .B(N1025));
NOR2XL inst_cellmath__201_0_I674 (.Y(N1453), .A(N1027), .B(N1026));
NAND2XL inst_cellmath__201_0_I675 (.Y(N1454), .A(N1027), .B(N1026));
NOR2XL inst_cellmath__201_0_I676 (.Y(N1455), .A(N1029), .B(N1028));
NAND2XL inst_cellmath__201_0_I677 (.Y(N1456), .A(N1029), .B(N1028));
NOR2XL inst_cellmath__201_0_I678 (.Y(N1457), .A(N1031), .B(N1030));
NAND2XL inst_cellmath__201_0_I679 (.Y(N1458), .A(N1031), .B(N1030));
NOR2XL inst_cellmath__201_0_I680 (.Y(N1459), .A(N1033), .B(N1032));
NAND2XL inst_cellmath__201_0_I681 (.Y(N1460), .A(N1033), .B(N1032));
NOR2XL inst_cellmath__201_0_I682 (.Y(N1461), .A(N1035), .B(N1034));
NAND2XL inst_cellmath__201_0_I683 (.Y(N1462), .A(N1035), .B(N1034));
NOR2XL inst_cellmath__201_0_I684 (.Y(N1463), .A(N1037), .B(N1036));
NAND2XL inst_cellmath__201_0_I685 (.Y(N1464), .A(N1037), .B(N1036));
NOR2XL inst_cellmath__201_0_I686 (.Y(N1465), .A(N1039), .B(N1038));
NAND2XL inst_cellmath__201_0_I687 (.Y(N1466), .A(N1039), .B(N1038));
NOR2XL inst_cellmath__201_0_I688 (.Y(N1467), .A(N1040), .B(N1041));
NAND2XL inst_cellmath__201_0_I689 (.Y(N1468), .A(N1040), .B(N1041));
NOR2XL inst_cellmath__201_0_I690 (.Y(N1469), .A(N1042), .B(N1043));
NAND2XL inst_cellmath__201_0_I691 (.Y(N1470), .A(N1042), .B(N1043));
NOR2XL inst_cellmath__201_0_I692 (.Y(N1471), .A(N1044), .B(N1045));
NAND2XL inst_cellmath__201_0_I693 (.Y(N1472), .A(N1044), .B(N1045));
NOR2XL inst_cellmath__201_0_I694 (.Y(N1473), .A(N1046), .B(N1047));
NAND2XL inst_cellmath__201_0_I695 (.Y(N1474), .A(N1046), .B(N1047));
NOR2XL inst_cellmath__201_0_I696 (.Y(N1475), .A(N1049), .B(N1048));
NAND2XL inst_cellmath__201_0_I697 (.Y(N1476), .A(N1049), .B(N1048));
AOI21X4 inst_cellmath__201_0_I701 (.Y(N1480), .A0(N1416), .A1(N1413), .B0(N1415));
AOI21X2 inst_cellmath__201_0_I705 (.Y(N1484), .A0(N1420), .A1(N1417), .B0(N1419));
NAND2X2 inst_cellmath__201_0_I706 (.Y(N1485), .A(N1420), .B(N1418));
AOI21X4 inst_cellmath__201_0_I709 (.Y(N1488), .A0(N1424), .A1(N1421), .B0(N1423));
NAND2X4 inst_cellmath__201_0_I710 (.Y(N1489), .A(N1424), .B(N1422));
AOI21X4 inst_cellmath__201_0_I713 (.Y(N1492), .A0(N1428), .A1(N1425), .B0(N1427));
NAND2X4 inst_cellmath__201_0_I714 (.Y(N1493), .A(N1428), .B(N1426));
AOI21X4 inst_cellmath__201_0_I717 (.Y(N1496), .A0(N1432), .A1(N1429), .B0(N1431));
NAND2X4 inst_cellmath__201_0_I718 (.Y(N1497), .A(N1432), .B(N1430));
AOI21X4 inst_cellmath__201_0_I721 (.Y(N1500), .A0(N1436), .A1(N1433), .B0(N1435));
NAND2X4 inst_cellmath__201_0_I722 (.Y(N1501), .A(N1436), .B(N1434));
AOI21X1 inst_cellmath__201_0_I725 (.Y(N1504), .A0(N1440), .A1(N1437), .B0(N1439));
NAND2X2 inst_cellmath__201_0_I726 (.Y(N1505), .A(N1440), .B(N1438));
AOI21XL inst_cellmath__201_0_I729 (.Y(N1508), .A0(N1444), .A1(N1441), .B0(N1443));
NAND2X1 inst_cellmath__201_0_I730 (.Y(N1509), .A(N1444), .B(N1442));
AOI21XL inst_cellmath__201_0_I733 (.Y(N1512), .A0(N1448), .A1(N1445), .B0(N1447));
NAND2XL inst_cellmath__201_0_I734 (.Y(N1513), .A(N1448), .B(N1446));
AOI21XL inst_cellmath__201_0_I737 (.Y(N1516), .A0(N1452), .A1(N1449), .B0(N1451));
NAND2XL inst_cellmath__201_0_I738 (.Y(N1517), .A(N1452), .B(N1450));
INVXL inst_cellmath__201_0_I1372 (.Y(N2420), .A(N1454));
AOI21XL inst_cellmath__201_0_I741 (.Y(N1520), .A0(N1456), .A1(N1453), .B0(N1455));
NAND2XL inst_cellmath__201_0_I742 (.Y(N1521), .A(N1456), .B(N1454));
AOI21XL inst_cellmath__201_0_I753 (.Y(N1532), .A0(N1460), .A1(N1457), .B0(N1459));
NAND2XL inst_cellmath__201_0_I754 (.Y(N1533), .A(N1460), .B(N1458));
INVXL inst_cellmath__201_0_I1380 (.Y(N2428), .A(N1462));
AOI21XL inst_cellmath__201_0_I757 (.Y(N1536), .A0(N1464), .A1(N1461), .B0(N1463));
NAND2XL inst_cellmath__201_0_I758 (.Y(N1537), .A(N1464), .B(N1462));
AOI21XL inst_cellmath__201_0_I769 (.Y(N1548), .A0(N1468), .A1(N1465), .B0(N1467));
NAND2XL inst_cellmath__201_0_I770 (.Y(N1549), .A(N1468), .B(N1466));
INVXL inst_cellmath__201_0_I1388 (.Y(N2436), .A(N1470));
AOI21XL inst_cellmath__201_0_I773 (.Y(N1552), .A0(N1472), .A1(N1469), .B0(N1471));
NAND2XL inst_cellmath__201_0_I774 (.Y(N1553), .A(N1472), .B(N1470));
AOI21XL inst_cellmath__201_0_I785 (.Y(N1564), .A0(N1476), .A1(N1473), .B0(N1475));
NAND2XL inst_cellmath__201_0_I786 (.Y(N1565), .A(N1476), .B(N1474));
INVXL inst_cellmath__201_0_I1395 (.Y(N2443), .A(N1049));
NOR2XL inst_cellmath__201_0_I793 (.Y(N1572), .A(N2443), .B(N1564));
NOR2XL andori2bb1_A_I1574 (.Y(N2545), .A(N2420), .B(N1516));
NOR2XL andori2bb1_A_I1575 (.Y(N2452), .A(N2545), .B(N1453));
OA21X1 inst_cellmath__201_0_I1480 (.Y(N2454), .A0(N1521), .A1(N1516), .B0(N1520));
OR2XL inst_cellmath__201_0_I1481 (.Y(N2455), .A(N1521), .B(N1517));
NOR2XL andori2bb1_A_I1576 (.Y(N2552), .A(N2428), .B(N1532));
NOR2XL andori2bb1_A_I1577 (.Y(N2460), .A(N2552), .B(N1461));
OA21X1 inst_cellmath__201_0_I1484 (.Y(N2462), .A0(N1537), .A1(N1532), .B0(N1536));
OR2XL inst_cellmath__201_0_I1485 (.Y(N2463), .A(N1537), .B(N1533));
NOR2XL andori2bb1_A_I1578 (.Y(N2559), .A(N2436), .B(N1548));
NOR2XL andori2bb1_A_I1579 (.Y(N2468), .A(N2559), .B(N1469));
OA21X1 inst_cellmath__201_0_I1488 (.Y(N2470), .A0(N1553), .A1(N1548), .B0(N1552));
OR2XL inst_cellmath__201_0_I1489 (.Y(N2471), .A(N1553), .B(N1549));
OR2XL inst_cellmath__201_0_I1490 (.Y(N2477), .A(N2443), .B(N1565));
INVXL inst_cellmath__201_0_I1430 (.Y(N2478), .A(N1480));
OAI21X4 inst_cellmath__201_0_I827 (.Y(N1607), .A0(N1485), .A1(N1480), .B0(N1484));
OAI21X2 inst_cellmath__201_0_I829 (.Y(N1609), .A0(N1489), .A1(N1484), .B0(N1488));
NOR2XL inst_cellmath__201_0_I830 (.Y(N1610), .A(N1489), .B(N1485));
OAI21X4 inst_cellmath__201_0_I831 (.Y(N1611), .A0(N1493), .A1(N1488), .B0(N1492));
NOR2X4 inst_cellmath__201_0_I832 (.Y(N1612), .A(N1493), .B(N1489));
OAI21X1 inst_cellmath__201_0_I833 (.Y(N1613), .A0(N1497), .A1(N1492), .B0(N1496));
NOR2X2 inst_cellmath__201_0_I834 (.Y(N1614), .A(N1497), .B(N1493));
OAI21X4 inst_cellmath__201_0_I835 (.Y(N1615), .A0(N1501), .A1(N1496), .B0(N1500));
NOR2X4 inst_cellmath__201_0_I836 (.Y(N1616), .A(N1501), .B(N1497));
OAI21X1 inst_cellmath__201_0_I837 (.Y(N1617), .A0(N1505), .A1(N1500), .B0(N1504));
NOR2X2 inst_cellmath__201_0_I838 (.Y(N1618), .A(N1505), .B(N1501));
OAI21X1 inst_cellmath__201_0_I839 (.Y(N1619), .A0(N1509), .A1(N1504), .B0(N1508));
NOR2X1 inst_cellmath__201_0_I840 (.Y(N1620), .A(N1509), .B(N1505));
OAI21XL inst_cellmath__201_0_I841 (.Y(N1621), .A0(N1513), .A1(N1508), .B0(N1512));
NOR2XL inst_cellmath__201_0_I842 (.Y(N1622), .A(N1513), .B(N1509));
OAI21XL inst_cellmath__201_0_I843 (.Y(N1623), .A0(N2455), .A1(N1512), .B0(N2454));
NOR2XL inst_cellmath__201_0_I844 (.Y(N1624), .A(N2455), .B(N1513));
OAI21XL inst_cellmath__201_0_I845 (.Y(N1625), .A0(N2463), .A1(N2454), .B0(N2462));
NOR2XL inst_cellmath__201_0_I846 (.Y(N1626), .A(N2463), .B(N2455));
OAI21XL inst_cellmath__201_0_I847 (.Y(N1627), .A0(N2471), .A1(N2462), .B0(N2470));
NOR2XL inst_cellmath__201_0_I848 (.Y(N1628), .A(N2471), .B(N2463));
INVXL inst_cellmath__201_0_I1431 (.Y(N2479), .A(N2478));
INVXL inst_cellmath__201_0_I1432 (.Y(N2480), .A(N1607));
AOI21XL inst_cellmath__201_0_I853 (.Y(N1633), .A0(N1610), .A1(N2478), .B0(N1609));
AOI21X2 inst_cellmath__201_0_I855 (.Y(N1635), .A0(N1612), .A1(N1607), .B0(N1611));
AOI21X1 inst_cellmath__201_0_I857 (.Y(N1637), .A0(N1614), .A1(N1609), .B0(N1613));
NAND2X1 inst_cellmath__201_0_I858 (.Y(N1638), .A(N1614), .B(N1610));
AOI21X2 inst_cellmath__201_0_I859 (.Y(N1639), .A0(N1616), .A1(N1611), .B0(N1615));
NAND2XL inst_cellmath__201_0_I860 (.Y(N1640), .A(N1616), .B(N1612));
AOI21XL inst_cellmath__201_0_I861 (.Y(N1641), .A0(N1618), .A1(N1613), .B0(N1617));
NAND2XL inst_cellmath__201_0_I862 (.Y(N1642), .A(N1618), .B(N1614));
AOI21X2 inst_cellmath__201_0_I863 (.Y(N1643), .A0(N1620), .A1(N1615), .B0(N1619));
NAND2X1 inst_cellmath__201_0_I864 (.Y(N1644), .A(N1620), .B(N1616));
AOI21XL inst_cellmath__201_0_I865 (.Y(N1645), .A0(N1622), .A1(N1617), .B0(N1621));
NAND2XL inst_cellmath__201_0_I866 (.Y(N1646), .A(N1622), .B(N1618));
AOI21XL inst_cellmath__201_0_I867 (.Y(N1647), .A0(N1624), .A1(N1619), .B0(N1623));
NAND2XL inst_cellmath__201_0_I868 (.Y(N1648), .A(N1624), .B(N1620));
AOI21XL inst_cellmath__201_0_I869 (.Y(N1649), .A0(N1626), .A1(N1621), .B0(N1625));
NAND2XL inst_cellmath__201_0_I870 (.Y(N1650), .A(N1626), .B(N1622));
AOI21XL inst_cellmath__201_0_I871 (.Y(N1651), .A0(N1628), .A1(N1623), .B0(N1627));
NAND2XL inst_cellmath__201_0_I872 (.Y(N1652), .A(N1628), .B(N1624));
INVXL inst_cellmath__201_0_I1435 (.Y(N2483), .A(N2479));
INVXL inst_cellmath__201_0_I1436 (.Y(N2484), .A(N2480));
INVXL inst_cellmath__201_0_I1437 (.Y(N2485), .A(N1633));
INVX1 inst_cellmath__201_0_I1438 (.Y(N2486), .A(N1635));
OAI21X1 inst_cellmath__201_0_I889 (.Y(N1669), .A0(N1646), .A1(N1637), .B0(N1645));
NOR2X1 inst_cellmath__201_0_I890 (.Y(N1670), .A(N1646), .B(N1638));
OAI21X1 inst_cellmath__201_0_I891 (.Y(N1671), .A0(N1648), .A1(N1639), .B0(N1647));
NOR2XL inst_cellmath__201_0_I892 (.Y(N1672), .A(N1648), .B(N1640));
OAI21XL inst_cellmath__201_0_I893 (.Y(N1673), .A0(N1650), .A1(N1641), .B0(N1649));
NOR2XL inst_cellmath__201_0_I894 (.Y(N1674), .A(N1650), .B(N1642));
OAI21X2 inst_cellmath__201_0_I895 (.Y(N1675), .A0(N1652), .A1(N1643), .B0(N1651));
NOR2X1 inst_cellmath__201_0_I896 (.Y(N1676), .A(N1652), .B(N1644));
INVXL inst_cellmath__201_0_I1439 (.Y(N2487), .A(N2483));
INVXL inst_cellmath__201_0_I1440 (.Y(N2488), .A(N2484));
INVXL inst_cellmath__201_0_I1441 (.Y(N2489), .A(N2485));
INVXL inst_cellmath__201_0_I1442 (.Y(N2490), .A(N2486));
OA21X1 inst_cellmath__201_0_I1491 (.Y(N2491), .A0(N2479), .A1(N1638), .B0(N1637));
OA21X1 inst_cellmath__201_0_I2451 (.Y(N2492), .A0(N1640), .A1(N2480), .B0(N1639));
OA21X1 inst_cellmath__201_0_I1550 (.Y(N2493), .A0(N1642), .A1(N1633), .B0(N1641));
OA21X1 inst_cellmath__201_0_I1494 (.Y(N2494), .A0(N1644), .A1(N1635), .B0(N1643));
AOI21X2 inst_cellmath__201_0_I913 (.Y(N1693), .A0(N1670), .A1(N2483), .B0(N1669));
AOI21X2 inst_cellmath__201_0_I915 (.Y(N1695), .A0(N1672), .A1(N2484), .B0(N1671));
AOI21X1 inst_cellmath__201_0_I917 (.Y(N1697), .A0(N1674), .A1(N2485), .B0(N1673));
AOI21X2 inst_cellmath__201_0_I919 (.Y(N1699), .A0(N1676), .A1(N2486), .B0(N1675));
INVXL buf1_A_I2460 (.Y(N3749), .A(N1699));
INVXL buf1_A_I2461 (.Y(N2496), .A(N3749));
NAND2BXL inst_cellmath__201_0_I959 (.Y(N1739), .AN(N1415), .B(N1416));
NAND2BXL inst_cellmath__201_0_I962 (.Y(N1742), .AN(N1417), .B(N1418));
NAND2BXL inst_cellmath__201_0_I965 (.Y(N1745), .AN(N1419), .B(N1420));
NAND2BXL inst_cellmath__201_0_I968 (.Y(N1748), .AN(N1421), .B(N1422));
NAND2BXL inst_cellmath__201_0_I971 (.Y(N1751), .AN(N1423), .B(N1424));
NAND2BXL inst_cellmath__201_0_I974 (.Y(N1754), .AN(N1425), .B(N1426));
NAND2BXL inst_cellmath__201_0_I977 (.Y(N1757), .AN(N1427), .B(N1428));
NAND2BXL inst_cellmath__201_0_I980 (.Y(N1760), .AN(N1429), .B(N1430));
NAND2BXL inst_cellmath__201_0_I983 (.Y(N1763), .AN(N1431), .B(N1432));
NAND2BXL inst_cellmath__201_0_I986 (.Y(N1766), .AN(N1433), .B(N1434));
NAND2BXL inst_cellmath__201_0_I989 (.Y(N1769), .AN(N1435), .B(N1436));
NAND2BXL inst_cellmath__201_0_I992 (.Y(N1772), .AN(N1437), .B(N1438));
NAND2BXL inst_cellmath__201_0_I995 (.Y(N1775), .AN(N1439), .B(N1440));
NAND2BXL inst_cellmath__201_0_I998 (.Y(N1778), .AN(N1441), .B(N1442));
NAND2BXL inst_cellmath__201_0_I1001 (.Y(N1781), .AN(N1443), .B(N1444));
NAND2BXL inst_cellmath__201_0_I1004 (.Y(N1784), .AN(N1445), .B(N1446));
NAND2BXL inst_cellmath__201_0_I1007 (.Y(N1787), .AN(N1447), .B(N1448));
NAND2BXL inst_cellmath__201_0_I1010 (.Y(N1790), .AN(N1449), .B(N1450));
NAND2BXL inst_cellmath__201_0_I1013 (.Y(N1793), .AN(N1451), .B(N1452));
NAND2BXL inst_cellmath__201_0_I1016 (.Y(N2058), .AN(N1453), .B(N1454));
NAND2BXL inst_cellmath__201_0_I1019 (.Y(N2069), .AN(N1455), .B(N1456));
NAND2BXL inst_cellmath__201_0_I1022 (.Y(N1802), .AN(N1457), .B(N1458));
NAND2BXL inst_cellmath__201_0_I1025 (.Y(N1805), .AN(N1459), .B(N1460));
NAND2BXL inst_cellmath__201_0_I1028 (.Y(N2087), .AN(N1461), .B(N1462));
NAND2BXL inst_cellmath__201_0_I1031 (.Y(N2098), .AN(N1463), .B(N1464));
NAND2BXL inst_cellmath__201_0_I1034 (.Y(N1814), .AN(N1465), .B(N1466));
NAND2BXL inst_cellmath__201_0_I1037 (.Y(N1817), .AN(N1467), .B(N1468));
NAND2BXL inst_cellmath__201_0_I1040 (.Y(N2116), .AN(N1469), .B(N1470));
NAND2BXL inst_cellmath__201_0_I1043 (.Y(N2127), .AN(N1471), .B(N1472));
NAND2BXL inst_cellmath__201_0_I1046 (.Y(N1826), .AN(N1473), .B(N1474));
NAND2BXL inst_cellmath__201_0_I1049 (.Y(N1829), .AN(N1475), .B(N1476));
XOR2XL inst_cellmath__201_0_I1495 (.Y(inst_cellmath__201_0_out0[17]), .A(N1413), .B(N1739));
XNOR2X1 inst_cellmath__201_0_I1055 (.Y(inst_cellmath__201_0_out0[18]), .A(N2487), .B(N1742));
XNOR2X1 inst_cellmath__201_0_I1056 (.Y(inst_cellmath__201_0_out0[20]), .A(N2488), .B(N1748));
XNOR2X1 inst_cellmath__201_0_I1057 (.Y(inst_cellmath__201_0_out0[22]), .A(N2489), .B(N1754));
XNOR2X1 inst_cellmath__201_0_I1058 (.Y(inst_cellmath__201_0_out0[24]), .A(N2490), .B(N1760));
XNOR2X1 inst_cellmath__201_0_I1059 (.Y(inst_cellmath__201_0_out0[26]), .A(N2491), .B(N1766));
XNOR2X1 inst_cellmath__201_0_I1060 (.Y(inst_cellmath__201_0_out0[28]), .A(N2492), .B(N1772));
XNOR2X1 inst_cellmath__201_0_I1061 (.Y(inst_cellmath__201_0_out0[30]), .A(N2493), .B(N1778));
XNOR2X1 inst_cellmath__201_0_I1062 (.Y(inst_cellmath__201_0_out0[32]), .A(N2494), .B(N1784));
XNOR2X1 inst_cellmath__201_0_I1063 (.Y(inst_cellmath__201_0_out0[34]), .A(N1693), .B(N1790));
XNOR2XL inst_cellmath__201_0_I2452 (.Y(inst_cellmath__201_0_out0[38]), .A(N1695), .B(N1802));
XNOR2X1 inst_cellmath__201_0_I1065 (.Y(inst_cellmath__201_0_out0[42]), .A(N1697), .B(N1814));
XNOR2XL inst_cellmath__201_0_I2453 (.Y(inst_cellmath__201_0_out0[46]), .A(N2496), .B(N1826));
XOR2XL node_cs_reduced_ii_local_A_I1496 (.Y(N1849), .A(N1745), .B(N1418));
XOR2XL node_cs_reduced_ii_local_A_I1497 (.Y(N1848), .A(N1745), .B(N1417));
MX2XL inst_cellmath__201_0_I1068 (.Y(inst_cellmath__201_0_out0[19]), .A(N1849), .B(N1848), .S0(N2487));
XOR2XL node_cs_reduced_ii_local_A_I1498 (.Y(N1852), .A(N1751), .B(N1422));
XOR2XL node_cs_reduced_ii_local_A_I1499 (.Y(N1851), .A(N1421), .B(N1751));
MX2XL inst_cellmath__201_0_I1070 (.Y(inst_cellmath__201_0_out0[21]), .A(N1852), .B(N1851), .S0(N2488));
XOR2XL node_cs_reduced_ii_local_A_I1500 (.Y(N1855), .A(N1426), .B(N1757));
XOR2XL node_cs_reduced_ii_local_A_I1501 (.Y(N1854), .A(N1425), .B(N1757));
MX2XL inst_cellmath__201_0_I1072 (.Y(inst_cellmath__201_0_out0[23]), .A(N1855), .B(N1854), .S0(N2489));
XOR2XL node_cs_reduced_ii_local_A_I1502 (.Y(N1858), .A(N1763), .B(N1430));
XOR2XL node_cs_reduced_ii_local_A_I1503 (.Y(N1857), .A(N1429), .B(N1763));
MX2XL inst_cellmath__201_0_I1074 (.Y(inst_cellmath__201_0_out0[25]), .A(N1858), .B(N1857), .S0(N2490));
XOR2XL node_cs_reduced_ii_local_A_I1504 (.Y(N1861), .A(N1434), .B(N1769));
XOR2XL node_cs_reduced_ii_local_A_I1505 (.Y(N1860), .A(N1769), .B(N1433));
MX2XL inst_cellmath__201_0_I1076 (.Y(inst_cellmath__201_0_out0[27]), .A(N1861), .B(N1860), .S0(N2491));
XOR2XL node_cs_reduced_ii_local_A_I1506 (.Y(N1864), .A(N1775), .B(N1438));
XOR2XL node_cs_reduced_ii_local_A_I1507 (.Y(N1863), .A(N1775), .B(N1437));
MX2XL inst_cellmath__201_0_I1078 (.Y(inst_cellmath__201_0_out0[29]), .A(N1864), .B(N1863), .S0(N2492));
XOR2XL node_cs_reduced_ii_local_A_I1508 (.Y(N1867), .A(N1781), .B(N1442));
XOR2XL node_cs_reduced_ii_local_A_I1509 (.Y(N1866), .A(N1781), .B(N1441));
MX2XL inst_cellmath__201_0_I1080 (.Y(inst_cellmath__201_0_out0[31]), .A(N1867), .B(N1866), .S0(N2493));
XOR2XL node_cs_reduced_ii_local_A_I1510 (.Y(N1870), .A(N1787), .B(N1446));
XOR2XL node_cs_reduced_ii_local_A_I1511 (.Y(N1869), .A(N1787), .B(N1445));
MX2XL inst_cellmath__201_0_I1082 (.Y(inst_cellmath__201_0_out0[33]), .A(N1870), .B(N1869), .S0(N2494));
XOR2XL node_cs_reduced_ii_local_A_I1512 (.Y(N1873), .A(N1793), .B(N1450));
XOR2XL node_cs_reduced_ii_local_A_I1513 (.Y(N1872), .A(N1793), .B(N1449));
MX2XL inst_cellmath__201_0_I1084 (.Y(inst_cellmath__201_0_out0[35]), .A(N1873), .B(N1872), .S0(N1693));
XOR2XL node_cs_ii_local_alt_A_I1163 (.Y(N1875), .A(N2058), .B(N1516));
NAND2XL node_cs_ii_local_alt_A_I1164 (.Y(N2056), .A(N1517), .B(N1516));
XNOR2X1 node_cs_ii_local_alt_A_I1165 (.Y(N1876), .A(N2058), .B(N2056));
MXI2XL inst_cellmath__201_0_I1086 (.Y(inst_cellmath__201_0_out0[36]), .A(N1876), .B(N1875), .S0(N1693));
XOR2XL node_cs_ii_local_alt_A_I1167 (.Y(N1878), .A(N2069), .B(N2452));
OAI21XL node_cs_ii_local_alt_A_I1514 (.Y(N2067), .A0(N2420), .A1(N1517), .B0(N2452));
XNOR2X1 node_cs_ii_local_alt_A_I1169 (.Y(N1879), .A(N2069), .B(N2067));
MXI2XL inst_cellmath__201_0_I1088 (.Y(inst_cellmath__201_0_out0[37]), .A(N1879), .B(N1878), .S0(N1693));
XOR2XL node_cs_reduced_ii_local_A_I1515 (.Y(N1882), .A(N1805), .B(N1458));
XOR2XL node_cs_reduced_ii_local_A_I1516 (.Y(N1881), .A(N1805), .B(N1457));
MX2XL inst_cellmath__201_0_I1090 (.Y(inst_cellmath__201_0_out0[39]), .A(N1882), .B(N1881), .S0(N1695));
XOR2XL node_cs_ii_local_alt_A_I1173 (.Y(N1884), .A(N2087), .B(N1532));
NAND2XL node_cs_ii_local_alt_A_I1174 (.Y(N2085), .A(N1533), .B(N1532));
XNOR2X1 node_cs_ii_local_alt_A_I1175 (.Y(N1885), .A(N2087), .B(N2085));
MXI2XL inst_cellmath__201_0_I1092 (.Y(inst_cellmath__201_0_out0[40]), .A(N1885), .B(N1884), .S0(N1695));
XOR2XL node_cs_ii_local_alt_A_I1177 (.Y(N1887), .A(N2098), .B(N2460));
OAI21XL node_cs_ii_local_alt_A_I1517 (.Y(N2096), .A0(N2428), .A1(N1533), .B0(N2460));
XNOR2X1 node_cs_ii_local_alt_A_I1179 (.Y(N1888), .A(N2098), .B(N2096));
MXI2XL inst_cellmath__201_0_I1094 (.Y(inst_cellmath__201_0_out0[41]), .A(N1888), .B(N1887), .S0(N1695));
XOR2XL node_cs_reduced_ii_local_A_I1518 (.Y(N1891), .A(N1817), .B(N1466));
XOR2XL node_cs_reduced_ii_local_A_I1519 (.Y(N1890), .A(N1817), .B(N1465));
MX2XL inst_cellmath__201_0_I1096 (.Y(inst_cellmath__201_0_out0[43]), .A(N1891), .B(N1890), .S0(N1697));
XOR2XL node_cs_ii_local_alt_A_I1183 (.Y(N1893), .A(N2116), .B(N1548));
NAND2XL node_cs_ii_local_alt_A_I1184 (.Y(N2114), .A(N1549), .B(N1548));
XNOR2X1 node_cs_ii_local_alt_A_I1185 (.Y(N1894), .A(N2116), .B(N2114));
MXI2XL inst_cellmath__201_0_I1098 (.Y(inst_cellmath__201_0_out0[44]), .A(N1894), .B(N1893), .S0(N1697));
XOR2XL node_cs_ii_local_alt_A_I1187 (.Y(N1896), .A(N2127), .B(N2468));
OAI21XL node_cs_ii_local_alt_A_I1520 (.Y(N2125), .A0(N2436), .A1(N1549), .B0(N2468));
XNOR2X1 node_cs_ii_local_alt_A_I1189 (.Y(N1897), .A(N2127), .B(N2125));
MXI2XL inst_cellmath__201_0_I1100 (.Y(inst_cellmath__201_0_out0[45]), .A(N1897), .B(N1896), .S0(N1697));
XOR2XL node_cs_reduced_ii_local_A_I1521 (.Y(N1900), .A(N1829), .B(N1474));
XOR2XL node_cs_reduced_ii_local_A_I1522 (.Y(N1899), .A(N1829), .B(N1473));
MX2XL inst_cellmath__201_0_I1102 (.Y(inst_cellmath__201_0_out0[47]), .A(N1900), .B(N1899), .S0(N2496));
XOR2XL node_cs_ii_local_alt_A_I1193 (.Y(N1902), .A(N2443), .B(N1564));
NAND2XL node_cs_ii_local_alt_A_I1194 (.Y(N2143), .A(N1565), .B(N1564));
XNOR2X1 node_cs_ii_local_alt_A_I1195 (.Y(N1903), .A(N2443), .B(N2143));
MXI2XL inst_cellmath__201_0_I1104 (.Y(inst_cellmath__201_0_out0[48]), .A(N1903), .B(N1902), .S0(N2496));
AOI2BB1X1 inst_cellmath__201_0_I1450 (.Y(N1907), .A0N(N2477), .A1N(N1699), .B0(N1572));
INVX1 inst_cellmath__201_0_I1449 (.Y(inst_cellmath__201_0_out0[49]), .A(N1907));
assign inst_cellmath__203__W1[0] = inst_cellmath__201_0_in1[0];
assign inst_cellmath__203__W1[1] = inst_cellmath__201_0_in0[1];
assign inst_cellmath__203__W1[2] = inst_cellmath__201_0_in0[2];
assign inst_cellmath__203__W1[3] = inst_cellmath__201_0_in0[3];
assign inst_cellmath__203__W1[4] = inst_cellmath__201_0_in0[4];
assign inst_cellmath__203__W1[5] = inst_cellmath__201_0_in0[5];
assign inst_cellmath__203__W1[6] = inst_cellmath__201_0_in0[6];
assign inst_cellmath__203__W1[7] = inst_cellmath__201_0_in0[7];
assign inst_cellmath__203__W1[8] = inst_cellmath__201_0_in0[8];
assign inst_cellmath__203__W1[9] = inst_cellmath__201_0_in0[9];
assign inst_cellmath__203__W1[10] = inst_cellmath__201_0_in0[10];
assign inst_cellmath__203__W1[11] = inst_cellmath__201_0_in0[11];
assign inst_cellmath__203__W1[12] = inst_cellmath__201_0_in0[12];
assign inst_cellmath__203__W1[13] = inst_cellmath__201_0_in0[13];
assign inst_cellmath__203__W1[14] = inst_cellmath__201_0_in0[14];
assign inst_cellmath__203__W1[15] = inst_cellmath__201_0_in0[15];
assign inst_cellmath__203__W1[16] = inst_cellmath__201_0_in0[16];
assign inst_cellmath__203__W1[17] = inst_cellmath__201_0_in0[17];
assign inst_cellmath__203__W1[18] = inst_cellmath__201_0_in0[18];
assign inst_cellmath__203__W1[19] = inst_cellmath__201_0_in0[19];
assign inst_cellmath__203__W1[20] = inst_cellmath__201_0_in0[20];
assign inst_cellmath__203__W1[21] = inst_cellmath__201_0_in0[21];
assign inst_cellmath__203__W1[22] = inst_cellmath__201_0_in0[22];
assign inst_cellmath__203__W1[23] = inst_cellmath__201_0_in0[23];
assign inst_cellmath__203__W1[24] = inst_cellmath__201_0_in0[24];
assign inst_cellmath__203__W1[25] = inst_cellmath__201_0_in0[25];
assign inst_cellmath__203__W1[26] = inst_cellmath__201_0_in0[26];
assign inst_cellmath__203__W1[27] = inst_cellmath__201_0_in0[27];
assign inst_cellmath__203__W1[28] = inst_cellmath__201_0_in0[28];
assign inst_cellmath__203__W1[29] = inst_cellmath__201_0_in0[29];
assign inst_cellmath__203__W1[30] = inst_cellmath__201_0_in0[30];
assign inst_cellmath__203__W1[31] = inst_cellmath__201_0_in0[31];
assign inst_cellmath__203__W1[32] = inst_cellmath__201_0_in1[32];
assign inst_cellmath__203__W1[33] = inst_cellmath__201_0_in1[33];
assign inst_cellmath__203__W1[34] = inst_cellmath__201_0_in0[34];
assign inst_cellmath__203__W1[35] = inst_cellmath__201_0_in1[35];
assign inst_cellmath__203__W1[36] = inst_cellmath__201_0_in0[36];
assign inst_cellmath__203__W1[37] = inst_cellmath__201_0_in0[37];
assign inst_cellmath__203__W1[38] = inst_cellmath__201_0_in0[38];
assign inst_cellmath__203__W1[39] = inst_cellmath__201_0_in0[39];
assign inst_cellmath__203__W1[40] = inst_cellmath__201_0_in0[40];
assign inst_cellmath__203__W1[41] = inst_cellmath__201_0_in0[41];
assign inst_cellmath__203__W1[42] = inst_cellmath__201_0_in0[42];
assign inst_cellmath__203__W1[43] = inst_cellmath__201_0_in0[43];
assign inst_cellmath__203__W1[44] = inst_cellmath__201_0_in0[44];
assign inst_cellmath__203__W1[45] = inst_cellmath__201_0_in0[45];
endmodule

module cynw_cm_float_sin_inst_cellmath__200_0_bdw1946085813_bdw (
	inst_cellmath__200_0_out0,
	inst_cellmath__200_0_in0
	); /* architecture "gate_level" */ 
output [48:0] inst_cellmath__200_0_out0;
input [49:0] inst_cellmath__200_0_in0;
wire N129,N130,N131,N132,N133,N134,N135 
	,N136,N137,N138,N139,N143,N145,N147,N148 
	,N252,N253,N254,N255,N256,N257,N258,N263 
	;
INVXL inst_cellmath__200_0_I28 (.Y(N129), .A(inst_cellmath__200_0_in0[28]));
INVXL inst_cellmath__200_0_I29 (.Y(N130), .A(inst_cellmath__200_0_in0[29]));
INVXL inst_cellmath__200_0_I30 (.Y(N131), .A(inst_cellmath__200_0_in0[30]));
INVXL inst_cellmath__200_0_I31 (.Y(N132), .A(inst_cellmath__200_0_in0[31]));
INVX1 inst_cellmath__200_0_I32 (.Y(N133), .A(inst_cellmath__200_0_in0[32]));
INVXL inst_cellmath__200_0_I33 (.Y(N134), .A(inst_cellmath__200_0_in0[33]));
INVXL inst_cellmath__200_0_I34 (.Y(N135), .A(inst_cellmath__200_0_in0[34]));
INVXL inst_cellmath__200_0_I35 (.Y(N136), .A(inst_cellmath__200_0_in0[35]));
INVXL inst_cellmath__200_0_I36 (.Y(N137), .A(inst_cellmath__200_0_in0[36]));
INVXL inst_cellmath__200_0_I37 (.Y(N138), .A(inst_cellmath__200_0_in0[37]));
INVXL inst_cellmath__200_0_I38 (.Y(N139), .A(inst_cellmath__200_0_in0[38]));
INVXL inst_cellmath__200_0_I42 (.Y(N143), .A(inst_cellmath__200_0_in0[42]));
INVXL inst_cellmath__200_0_I44 (.Y(N145), .A(inst_cellmath__200_0_in0[44]));
INVXL inst_cellmath__200_0_I46 (.Y(N147), .A(inst_cellmath__200_0_in0[46]));
INVXL inst_cellmath__200_0_I47 (.Y(N148), .A(inst_cellmath__200_0_in0[47]));
INVXL inst_cellmath__200_0_I107 (.Y(N258), .A(inst_cellmath__200_0_in0[49]));
CLKINVX4 inst_cellmath__200_0_I101 (.Y(N252), .A(inst_cellmath__200_0_in0[49]));
INVXL inst_cellmath__200_0_I112 (.Y(N263), .A(N258));
INVX2 inst_cellmath__200_0_I106 (.Y(N257), .A(N252));
CLKINVX4 inst_cellmath__200_0_I105 (.Y(N256), .A(N252));
INVX3 inst_cellmath__200_0_I104 (.Y(N255), .A(N252));
INVX3 inst_cellmath__200_0_I103 (.Y(N254), .A(N252));
INVX2 inst_cellmath__200_0_I102 (.Y(N253), .A(N252));
NOR2BX1 inst_cellmath__200_0_I786 (.Y(inst_cellmath__200_0_out0[0]), .AN(inst_cellmath__200_0_in0[0]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I787 (.Y(inst_cellmath__200_0_out0[1]), .AN(inst_cellmath__200_0_in0[1]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I788 (.Y(inst_cellmath__200_0_out0[2]), .AN(inst_cellmath__200_0_in0[2]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I789 (.Y(inst_cellmath__200_0_out0[3]), .AN(inst_cellmath__200_0_in0[3]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I790 (.Y(inst_cellmath__200_0_out0[4]), .AN(inst_cellmath__200_0_in0[4]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I791 (.Y(inst_cellmath__200_0_out0[5]), .AN(inst_cellmath__200_0_in0[5]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I792 (.Y(inst_cellmath__200_0_out0[6]), .AN(inst_cellmath__200_0_in0[6]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I793 (.Y(inst_cellmath__200_0_out0[7]), .AN(inst_cellmath__200_0_in0[7]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I794 (.Y(inst_cellmath__200_0_out0[8]), .AN(inst_cellmath__200_0_in0[8]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I795 (.Y(inst_cellmath__200_0_out0[9]), .AN(inst_cellmath__200_0_in0[9]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I796 (.Y(inst_cellmath__200_0_out0[10]), .AN(inst_cellmath__200_0_in0[10]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I797 (.Y(inst_cellmath__200_0_out0[11]), .AN(inst_cellmath__200_0_in0[11]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I798 (.Y(inst_cellmath__200_0_out0[12]), .AN(inst_cellmath__200_0_in0[12]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I799 (.Y(inst_cellmath__200_0_out0[13]), .AN(inst_cellmath__200_0_in0[13]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I800 (.Y(inst_cellmath__200_0_out0[14]), .AN(inst_cellmath__200_0_in0[14]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I801 (.Y(inst_cellmath__200_0_out0[15]), .AN(inst_cellmath__200_0_in0[15]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I802 (.Y(inst_cellmath__200_0_out0[16]), .AN(inst_cellmath__200_0_in0[16]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I803 (.Y(inst_cellmath__200_0_out0[17]), .AN(inst_cellmath__200_0_in0[17]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I804 (.Y(inst_cellmath__200_0_out0[18]), .AN(inst_cellmath__200_0_in0[18]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I805 (.Y(inst_cellmath__200_0_out0[19]), .AN(inst_cellmath__200_0_in0[19]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I806 (.Y(inst_cellmath__200_0_out0[20]), .AN(inst_cellmath__200_0_in0[20]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I807 (.Y(inst_cellmath__200_0_out0[21]), .AN(inst_cellmath__200_0_in0[21]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I808 (.Y(inst_cellmath__200_0_out0[22]), .AN(inst_cellmath__200_0_in0[22]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I809 (.Y(inst_cellmath__200_0_out0[23]), .AN(inst_cellmath__200_0_in0[23]), .B(N263));
NOR2BX1 inst_cellmath__200_0_I810 (.Y(inst_cellmath__200_0_out0[24]), .AN(inst_cellmath__200_0_in0[24]), .B(N257));
NOR2BX1 inst_cellmath__200_0_I811 (.Y(inst_cellmath__200_0_out0[25]), .AN(inst_cellmath__200_0_in0[25]), .B(N257));
NOR2BX1 inst_cellmath__200_0_I812 (.Y(inst_cellmath__200_0_out0[26]), .AN(inst_cellmath__200_0_in0[26]), .B(N257));
NOR2BX1 inst_cellmath__200_0_I813 (.Y(inst_cellmath__200_0_out0[27]), .AN(inst_cellmath__200_0_in0[27]), .B(N257));
NOR2X2 inst_cellmath__200_0_I77 (.Y(inst_cellmath__200_0_out0[28]), .A(N129), .B(N257));
NOR2X4 inst_cellmath__200_0_I78 (.Y(inst_cellmath__200_0_out0[29]), .A(N130), .B(N256));
NOR2X4 inst_cellmath__200_0_I79 (.Y(inst_cellmath__200_0_out0[30]), .A(N131), .B(N256));
NOR2X2 inst_cellmath__200_0_I80 (.Y(inst_cellmath__200_0_out0[31]), .A(N132), .B(N256));
NOR2X2 inst_cellmath__200_0_I81 (.Y(inst_cellmath__200_0_out0[32]), .A(N133), .B(N256));
NOR2X4 inst_cellmath__200_0_I82 (.Y(inst_cellmath__200_0_out0[33]), .A(N134), .B(N256));
NOR2X2 inst_cellmath__200_0_I83 (.Y(inst_cellmath__200_0_out0[34]), .A(N135), .B(N255));
NOR2X2 inst_cellmath__200_0_I84 (.Y(inst_cellmath__200_0_out0[35]), .A(N136), .B(N255));
NOR2X2 inst_cellmath__200_0_I85 (.Y(inst_cellmath__200_0_out0[36]), .A(N137), .B(N255));
NOR2X2 inst_cellmath__200_0_I86 (.Y(inst_cellmath__200_0_out0[37]), .A(N138), .B(N255));
NOR2X4 inst_cellmath__200_0_I87 (.Y(inst_cellmath__200_0_out0[38]), .A(N139), .B(N255));
NOR2BX2 inst_cellmath__200_0_I825 (.Y(inst_cellmath__200_0_out0[39]), .AN(inst_cellmath__200_0_in0[39]), .B(N254));
NOR2BX1 inst_cellmath__200_0_I826 (.Y(inst_cellmath__200_0_out0[40]), .AN(inst_cellmath__200_0_in0[40]), .B(N254));
NOR2BX1 inst_cellmath__200_0_I827 (.Y(inst_cellmath__200_0_out0[41]), .AN(inst_cellmath__200_0_in0[41]), .B(N254));
NOR2X2 inst_cellmath__200_0_I91 (.Y(inst_cellmath__200_0_out0[42]), .A(N143), .B(N254));
NOR2BX1 inst_cellmath__200_0_I829 (.Y(inst_cellmath__200_0_out0[43]), .AN(inst_cellmath__200_0_in0[43]), .B(N254));
NOR2X2 inst_cellmath__200_0_I93 (.Y(inst_cellmath__200_0_out0[44]), .A(N145), .B(N253));
NOR2BX2 inst_cellmath__200_0_I831 (.Y(inst_cellmath__200_0_out0[45]), .AN(inst_cellmath__200_0_in0[45]), .B(N253));
NOR2X4 inst_cellmath__200_0_I95 (.Y(inst_cellmath__200_0_out0[46]), .A(N147), .B(N253));
NOR2X2 inst_cellmath__200_0_I96 (.Y(inst_cellmath__200_0_out0[47]), .A(N148), .B(N253));
NOR2BX1 inst_cellmath__200_0_I834 (.Y(inst_cellmath__200_0_out0[48]), .AN(inst_cellmath__200_0_in0[48]), .B(N253));
endmodule

module cynw_cm_float_sin_inst_cellmath__19_0_bdw1946085813_bdw (
	inst_cellmath__19_0_out0,
	inst_cellmath__19_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19_0_out0;
input [7:0] inst_cellmath__19_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2X1 inst_cellmath__19_0_I0 (.Y(N11), .A(inst_cellmath__19_0_in0[7]), .B(inst_cellmath__19_0_in0[0]));
NAND2XL inst_cellmath__19_0_I1 (.Y(N12), .A(inst_cellmath__19_0_in0[6]), .B(inst_cellmath__19_0_in0[5]));
NAND2X1 inst_cellmath__19_0_I2 (.Y(N13), .A(inst_cellmath__19_0_in0[4]), .B(inst_cellmath__19_0_in0[3]));
NAND2XL inst_cellmath__19_0_I3 (.Y(N14), .A(inst_cellmath__19_0_in0[2]), .B(inst_cellmath__19_0_in0[1]));
NOR2XL inst_cellmath__19_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__19_0_I5 (.Y(N16), .A(N13), .B(N14));
CLKAND2X2 inst_cellmath__19_0_I6 (.Y(inst_cellmath__19_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_sin_inst_cellmath__24_0_bdw1946085813_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48;
NOR2XL inst_cellmath__24_0_I0 (.Y(N26), .A(inst_cellmath__24_0_in0[0]), .B(inst_cellmath__24_0_in0[1]));
NOR2XL inst_cellmath__24_0_I1 (.Y(N27), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
NOR2XL inst_cellmath__24_0_I2 (.Y(N28), .A(inst_cellmath__24_0_in0[20]), .B(inst_cellmath__24_0_in0[19]));
NOR2XL inst_cellmath__24_0_I3 (.Y(N29), .A(inst_cellmath__24_0_in0[18]), .B(inst_cellmath__24_0_in0[17]));
NOR2XL inst_cellmath__24_0_I4 (.Y(N30), .A(inst_cellmath__24_0_in0[16]), .B(inst_cellmath__24_0_in0[15]));
NOR2XL inst_cellmath__24_0_I5 (.Y(N31), .A(inst_cellmath__24_0_in0[14]), .B(inst_cellmath__24_0_in0[13]));
NOR2XL inst_cellmath__24_0_I6 (.Y(N32), .A(inst_cellmath__24_0_in0[12]), .B(inst_cellmath__24_0_in0[11]));
NOR2XL inst_cellmath__24_0_I7 (.Y(N33), .A(inst_cellmath__24_0_in0[10]), .B(inst_cellmath__24_0_in0[9]));
NOR2XL inst_cellmath__24_0_I8 (.Y(N34), .A(inst_cellmath__24_0_in0[8]), .B(inst_cellmath__24_0_in0[7]));
NOR2XL inst_cellmath__24_0_I9 (.Y(N35), .A(inst_cellmath__24_0_in0[6]), .B(inst_cellmath__24_0_in0[5]));
NOR2XL inst_cellmath__24_0_I10 (.Y(N36), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in0[3]));
INVXL inst_cellmath__24_0_I11 (.Y(N37), .A(inst_cellmath__24_0_in0[2]));
NAND2XL inst_cellmath__24_0_I12 (.Y(N38), .A(N37), .B(N26));
NAND2XL inst_cellmath__24_0_I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__24_0_I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__24_0_I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__24_0_I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__24_0_I17 (.Y(N43), .A(N35), .B(N36));
NOR2XL inst_cellmath__24_0_I18 (.Y(N44), .A(N38), .B(N39));
NOR2XL inst_cellmath__24_0_I19 (.Y(N45), .A(N40), .B(N41));
NAND2XL inst_cellmath__24_0_I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__24_0_I169 (.Y(N48), .A(N42), .B(N43));
NOR2XL inst_cellmath__24_0_I23 (.Y(inst_cellmath__24_0_out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_sin_inst_cellmath__66_0_bdw1946085813_bdw (
	inst_cellmath__66_0_out0,
	inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__66_0_out0;
input  inst_cellmath__66_0_in0,
	inst_cellmath__66_0_in1,
	inst_cellmath__66_0_in2;
wire N6,N8;
INVXL inst_cellmath__66_0_I0 (.Y(N6), .A(inst_cellmath__66_0_in2));
CLKAND2X3 inst_cellmath__66_0_I1 (.Y(N8), .A(N6), .B(inst_cellmath__66_0_in1));
CLKAND2X3 inst_cellmath__66_0_I3 (.Y(inst_cellmath__66_0_out0), .A(N8), .B(inst_cellmath__66_0_in0));
endmodule

module cynw_cm_float_sin_inst_cellmath__67_0_bdw1946085813_bdw (
	inst_cellmath__67_0_out0,
	inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__67_0_out0;
input  inst_cellmath__67_0_in0,
	inst_cellmath__67_0_in1,
	inst_cellmath__67_0_in2;
wire N7;
CLKAND2X2 inst_cellmath__67_0_I0 (.Y(N7), .A(inst_cellmath__67_0_in2), .B(inst_cellmath__67_0_in1));
CLKAND2X3 inst_cellmath__67_0_I2 (.Y(inst_cellmath__67_0_out0), .A(N7), .B(inst_cellmath__67_0_in0));
endmodule

module cynw_cm_float_sin_inst_cellmath__68_0_bdw1946085813_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__68_0_out0;
input  inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1;
OR2XL inst_cellmath__68_0_I0 (.Y(inst_cellmath__68_0_out0), .A(inst_cellmath__68_0_in0), .B(inst_cellmath__68_0_in1));
endmodule

module cynw_cm_float_sin_inst_cellmath__69_0_bdw1946085813_bdw (
	inst_cellmath__69_0_out0,
	inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__69_0_out0;
input  inst_cellmath__69_0_in0,
	inst_cellmath__69_0_in1;
wire N5;
INVXL inst_cellmath__69_0_I0 (.Y(N5), .A(inst_cellmath__69_0_in1));
NOR2X2 inst_cellmath__69_0_I1 (.Y(inst_cellmath__69_0_out0), .A(N5), .B(inst_cellmath__69_0_in0));
endmodule

module cynw_cm_float_sin_inst_cellmath__82_0_bdw1946085813_bdw (
	inst_cellmath__82_0_out0,
	inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__82_0_out0;
input  inst_cellmath__82_0_in0,
	inst_cellmath__82_0_in1;
wire N5;
NOR2XL inst_cellmath__82_0_I0 (.Y(N5), .A(inst_cellmath__82_0_in1), .B(inst_cellmath__82_0_in0));
INVXL inst_cellmath__82_0_I1 (.Y(inst_cellmath__82_0_out0), .A(N5));
endmodule

module cynw_cm_float_sin_inst_cellmath__17_0_bdw1946085813_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NOR2X1 inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[0]));
NOR2X1 inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[6]), .B(inst_cellmath__17_0_in0[5]));
NOR2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[4]), .B(inst_cellmath__17_0_in0[3]));
NOR2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[2]), .B(inst_cellmath__17_0_in0[1]));
NAND2X1 inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_sin_inst_cellmath__79__46__bdw1946085813_bdw (
	inst_cellmath__79__46__out0,
	inst_cellmath__79__46__in0,
	inst_cellmath__79__46__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__79__46__out0;
input  inst_cellmath__79__46__in0,
	inst_cellmath__79__46__in1;
OR2XL inst_cellmath__79__46__I0 (.Y(inst_cellmath__79__46__out0[0]), .A(inst_cellmath__79__46__in1), .B(inst_cellmath__79__46__in0));
endmodule

module cynw_cm_float_sin_inst_cellmath__228__231__bdw1946085813_bdw (
	inst_cellmath__228__231__out0,
	inst_cellmath__228__231__in0,
	inst_cellmath__228__231__in1,
	inst_cellmath__228__231__in2
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__228__231__out0;
input  inst_cellmath__228__231__in0;
input [0:0] inst_cellmath__228__231__in1;
input  inst_cellmath__228__231__in2;
OR3XL inst_cellmath__228__231__I4 (.Y(inst_cellmath__228__231__out0[0]), .A(inst_cellmath__228__231__in0), .B(inst_cellmath__228__231__in2), .C(inst_cellmath__228__231__in1[0]));
endmodule

module cynw_cm_float_sin_inst_cellmath__216__184__bdw1946085813_bdw (
	inst_cellmath__216__184__out0,
	inst_cellmath__216__184__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__216__184__out0;
input [7:0] inst_cellmath__216__184__in0;
wire N56,N58,N60;
NAND2X1 inst_cellmath__216__184__I31 (.Y(N56), .A(inst_cellmath__216__184__in0[4]), .B(inst_cellmath__216__184__in0[3]));
NAND2X1 inst_cellmath__216__184__I32 (.Y(N58), .A(inst_cellmath__216__184__in0[5]), .B(inst_cellmath__216__184__in0[6]));
NOR2X1 inst_cellmath__216__184__I33 (.Y(N60), .A(N56), .B(N58));
NOR2X1 inst_cellmath__216__184__I34 (.Y(inst_cellmath__216__184__out0[0]), .A(inst_cellmath__216__184__in0[7]), .B(N60));
endmodule

module cynw_cm_float_sin_inst_cellmath__219_0_bdw1946085813_bdw (
	inst_cellmath__219_0_out0,
	inst_cellmath__219_0_in0,
	inst_cellmath__219_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__219_0_out0;
input [22:22] inst_cellmath__219_0_in0;
input [48:48] inst_cellmath__219_0_in1;
AND2XL inst_cellmath__219_0_I0 (.Y(inst_cellmath__219_0_out0), .A(inst_cellmath__219_0_in0[22]), .B(inst_cellmath__219_0_in1[48]));
endmodule

module cynw_cm_float_sin_inst_cellmath__211__182__bdw1946085813_bdw (
	inst_cellmath__211__182__out0,
	inst_cellmath__211__182__in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__211__182__out0;
input [47:25] inst_cellmath__211__182__in0;
wire N100,N106,N108,N109,N112,N113,N114 
	,N115,N116,N117,N118,N119,N120,N121,N122 
	,N123,N124,N125,N126,N127,N128,N129,N131 
	,N132,N133,N135,N136,N137,N139,N140,N141 
	,N155,N157,N158,N160,N162,N163,N164,N165 
	,N166,N167,N168,N171,N172,N180,N182,N183 
	,N189,N191,N194,N216,N218,N232,N234,N236 
	,N240,N242,N282;
INVX1 inst_cellmath__211__182__I7 (.Y(N100), .A(inst_cellmath__211__182__in0[47]));
INVXL inst_cellmath__211__182__I11 (.Y(N106), .A(inst_cellmath__211__182__in0[25]));
INVXL inst_cellmath__211__182__I12 (.Y(N108), .A(inst_cellmath__211__182__in0[27]));
OAI21X2 inst_cellmath__211__182__I13 (.Y(N109), .A0(inst_cellmath__211__182__in0[26]), .A1(N106), .B0(N108));
OR2XL inst_cellmath__211__182__I15 (.Y(N155), .A(inst_cellmath__211__182__in0[27]), .B(inst_cellmath__211__182__in0[26]));
INVX1 inst_cellmath__211__182__I16 (.Y(N112), .A(inst_cellmath__211__182__in0[28]));
NOR2X2 inst_cellmath__211__182__I17 (.Y(N113), .A(inst_cellmath__211__182__in0[29]), .B(N112));
INVX1 inst_cellmath__211__182__I18 (.Y(N114), .A(inst_cellmath__211__182__in0[31]));
OAI21X4 inst_cellmath__211__182__I19 (.Y(N115), .A0(inst_cellmath__211__182__in0[30]), .A1(N113), .B0(N114));
NOR2X4 inst_cellmath__211__182__I20 (.Y(N116), .A(inst_cellmath__211__182__in0[29]), .B(inst_cellmath__211__182__in0[28]));
NOR2X4 inst_cellmath__211__182__I21 (.Y(N117), .A(inst_cellmath__211__182__in0[31]), .B(inst_cellmath__211__182__in0[30]));
INVX1 inst_cellmath__211__182__I22 (.Y(N118), .A(inst_cellmath__211__182__in0[32]));
NOR2X2 inst_cellmath__211__182__I23 (.Y(N119), .A(inst_cellmath__211__182__in0[33]), .B(N118));
INVX1 inst_cellmath__211__182__I24 (.Y(N120), .A(inst_cellmath__211__182__in0[35]));
OAI21X2 inst_cellmath__211__182__I25 (.Y(N121), .A0(inst_cellmath__211__182__in0[34]), .A1(N119), .B0(N120));
NOR2X4 inst_cellmath__211__182__I26 (.Y(N122), .A(inst_cellmath__211__182__in0[33]), .B(inst_cellmath__211__182__in0[32]));
NOR2X4 inst_cellmath__211__182__I27 (.Y(N123), .A(inst_cellmath__211__182__in0[35]), .B(inst_cellmath__211__182__in0[34]));
INVX1 inst_cellmath__211__182__I28 (.Y(N124), .A(inst_cellmath__211__182__in0[36]));
NOR2X2 inst_cellmath__211__182__I29 (.Y(N125), .A(inst_cellmath__211__182__in0[37]), .B(N124));
INVX1 inst_cellmath__211__182__I30 (.Y(N126), .A(inst_cellmath__211__182__in0[39]));
OAI21X4 inst_cellmath__211__182__I31 (.Y(N127), .A0(inst_cellmath__211__182__in0[38]), .A1(N125), .B0(N126));
NOR2X4 inst_cellmath__211__182__I32 (.Y(N128), .A(inst_cellmath__211__182__in0[37]), .B(inst_cellmath__211__182__in0[36]));
NOR2X6 inst_cellmath__211__182__I33 (.Y(N129), .A(inst_cellmath__211__182__in0[39]), .B(inst_cellmath__211__182__in0[38]));
NOR2BX1 inst_cellmath__211__182__I327 (.Y(N131), .AN(inst_cellmath__211__182__in0[40]), .B(inst_cellmath__211__182__in0[41]));
INVXL inst_cellmath__211__182__I36 (.Y(N132), .A(inst_cellmath__211__182__in0[43]));
OAI21X2 inst_cellmath__211__182__I37 (.Y(N133), .A0(inst_cellmath__211__182__in0[42]), .A1(N131), .B0(N132));
NOR2X1 inst_cellmath__211__182__I38 (.Y(N167), .A(inst_cellmath__211__182__in0[41]), .B(inst_cellmath__211__182__in0[40]));
NOR2X2 inst_cellmath__211__182__I39 (.Y(N135), .A(inst_cellmath__211__182__in0[43]), .B(inst_cellmath__211__182__in0[42]));
INVX2 inst_cellmath__211__182__I40 (.Y(N136), .A(inst_cellmath__211__182__in0[44]));
NOR2X2 inst_cellmath__211__182__I41 (.Y(N137), .A(inst_cellmath__211__182__in0[45]), .B(N136));
OAI21X4 inst_cellmath__211__182__I43 (.Y(N139), .A0(inst_cellmath__211__182__in0[46]), .A1(N137), .B0(N100));
NOR2X4 inst_cellmath__211__182__I44 (.Y(N140), .A(inst_cellmath__211__182__in0[45]), .B(inst_cellmath__211__182__in0[44]));
NOR2X4 inst_cellmath__211__182__I45 (.Y(N141), .A(inst_cellmath__211__182__in0[47]), .B(inst_cellmath__211__182__in0[46]));
INVXL inst_cellmath__211__182__I60 (.Y(N157), .A(N117));
AOI21XL inst_cellmath__211__182__I61 (.Y(N158), .A0(N116), .A1(N155), .B0(N157));
NAND2X2 inst_cellmath__211__182__I63 (.Y(N160), .A(N117), .B(N116));
NAND2BX1 inst_cellmath__211__182__I160 (.Y(N162), .AN(N122), .B(N123));
INVXL inst_cellmath__211__182__I66 (.Y(N163), .A(N129));
AOI21X1 inst_cellmath__211__182__I67 (.Y(N164), .A0(N128), .A1(N162), .B0(N163));
NAND2X4 inst_cellmath__211__182__I68 (.Y(N165), .A(N123), .B(N122));
NAND2X6 inst_cellmath__211__182__I69 (.Y(N166), .A(N129), .B(N128));
NAND2BXL inst_cellmath__211__182__I161 (.Y(N168), .AN(N167), .B(N135));
NAND2X2 inst_cellmath__211__182__I74 (.Y(N171), .A(N135), .B(N167));
NAND2X6 inst_cellmath__211__182__I75 (.Y(N172), .A(N141), .B(N140));
INVXL inst_cellmath__211__182__I83 (.Y(N180), .A(N160));
INVXL inst_cellmath__211__182__I84 (.Y(N182), .A(N166));
OAI21XL inst_cellmath__211__182__I85 (.Y(N183), .A0(N165), .A1(N180), .B0(N182));
NOR2X6 inst_cellmath__211__182__I87 (.Y(N194), .A(N166), .B(N165));
NAND2BXL inst_cellmath__211__182__I162 (.Y(N189), .AN(N172), .B(N171));
NOR2X4 inst_cellmath__211__182__I92 (.Y(N191), .A(N172), .B(N171));
NAND2BXL inst_cellmath__211__182__I186 (.Y(inst_cellmath__211__182__out0[3]), .AN(N194), .B(N191));
INVX3 inst_cellmath__211__182__I152 (.Y(N282), .A(N191));
INVXL inst_cellmath__211__182__I101 (.Y(inst_cellmath__211__182__out0[4]), .A(N282));
OAI21XL inst_cellmath__211__182__I106 (.Y(inst_cellmath__211__182__out0[2]), .A0(N282), .A1(N183), .B0(N189));
AOI21X2 inst_cellmath__211__182__I112 (.Y(N216), .A0(N194), .A1(N158), .B0(N164));
OAI2BB1X1 inst_cellmath__211__182__I172 (.Y(N218), .A0N(N140), .A1N(N168), .B0(N141));
OAI21X1 inst_cellmath__211__182__I116 (.Y(inst_cellmath__211__182__out0[1]), .A0(N282), .A1(N216), .B0(N218));
OAI21X4 inst_cellmath__211__182__I126 (.Y(N232), .A0(N160), .A1(N109), .B0(N115));
OAI21X4 inst_cellmath__211__182__I128 (.Y(N234), .A0(N166), .A1(N121), .B0(N127));
OAI21X2 inst_cellmath__211__182__I130 (.Y(N236), .A0(N172), .A1(N133), .B0(N139));
AOI21X4 inst_cellmath__211__182__I134 (.Y(N240), .A0(N194), .A1(N232), .B0(N234));
INVX2 inst_cellmath__211__182__I136 (.Y(N242), .A(N236));
OAI21X4 inst_cellmath__211__182__I138 (.Y(inst_cellmath__211__182__out0[0]), .A0(N282), .A1(N240), .B0(N242));
endmodule

module cynw_cm_float_sin_inst_cellmath__215_0_bdw1946085813_bdw (
	inst_cellmath__215_0_out0,
	inst_cellmath__215_0_in0
	); /* architecture "gate_level" */ 
output [4:0] inst_cellmath__215_0_out0;
input [4:0] inst_cellmath__215_0_in0;
wire N47,N67,N72,N89,N161,N171;
INVXL inst_cellmath__215_0_I85 (.Y(N161), .A(inst_cellmath__215_0_in0[0]));
AND2XL inst_cellmath__215_0_I21 (.Y(N47), .A(inst_cellmath__215_0_in0[1]), .B(inst_cellmath__215_0_in0[0]));
NAND2XL inst_cellmath__215_0_I24 (.Y(N89), .A(inst_cellmath__215_0_in0[2]), .B(inst_cellmath__215_0_in0[1]));
NOR2XL inst_cellmath__215_0_I33 (.Y(N67), .A(N89), .B(N161));
AO21XL inst_cellmath__215_0_I35 (.Y(N72), .A0(inst_cellmath__215_0_in0[2]), .A1(N47), .B0(inst_cellmath__215_0_in0[3]));
INVXL inst_cellmath__215_0_I64 (.Y(inst_cellmath__215_0_out0[0]), .A(inst_cellmath__215_0_in0[0]));
XNOR2X1 inst_cellmath__215_0_I100 (.Y(inst_cellmath__215_0_out0[1]), .A(N161), .B(inst_cellmath__215_0_in0[1]));
CLKXOR2X1 inst_cellmath__215_0_I130 (.Y(inst_cellmath__215_0_out0[2]), .A(N47), .B(inst_cellmath__215_0_in0[2]));
XNOR2X1 inst_cellmath__215_0_I98 (.Y(inst_cellmath__215_0_out0[3]), .A(N67), .B(inst_cellmath__215_0_in0[3]));
INVXL xnor2_A_I104 (.Y(N171), .A(N72));
MXI2XL xnor2_A_I105 (.Y(inst_cellmath__215_0_out0[4]), .A(N72), .B(N171), .S0(inst_cellmath__215_0_in0[4]));
endmodule

module cynw_cm_float_sin_inst_cellmath__220__188__bdw1946085813_bdw (
	inst_cellmath__220__188__out0,
	inst_cellmath__220__188__in0,
	inst_cellmath__220__188__in1
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__220__188__out0;
input [4:0] inst_cellmath__220__188__in0;
input [47:25] inst_cellmath__220__188__in1;
wire N55,N57,N58,N59,N60,N61,N62 
	,N63,N64,N65,N66,N67,N68,N69,N70 
	,N71,N72,N73,N74,N75,N76,N77,N78 
	,N106,N108,N110,N111,N112,N113,N114,N115 
	,N116,N117,N118,N119,N120,N121,N122,N123 
	,N124,N125,N126,N127,N128,N129,N130,N158 
	,N160,N162,N164,N166,N167,N168,N169,N170 
	,N171,N172,N173,N174,N175,N176,N177,N178 
	,N179,N180,N181,N182,N183,N184,N212,N214 
	,N216,N218,N220,N222,N224,N226,N228,N230 
	,N232,N234,N236,N238,N240,N242,N244,N245 
	,N246,N247,N248,N249,N250,N341,N342,N343 
	,N347,N348,N349,N351,N355,N357,N358,N360 
	,N364;
INVX2 inst_cellmath__220__188__I282 (.Y(N341), .A(inst_cellmath__220__188__in0[0]));
AND2XL inst_cellmath__220__188__I2 (.Y(N55), .A(N341), .B(inst_cellmath__220__188__in1[25]));
MX2XL inst_cellmath__220__188__I3 (.Y(N57), .A(inst_cellmath__220__188__in1[25]), .B(inst_cellmath__220__188__in1[26]), .S0(N341));
MX2XL inst_cellmath__220__188__I4 (.Y(N58), .A(inst_cellmath__220__188__in1[26]), .B(inst_cellmath__220__188__in1[27]), .S0(N341));
MX2XL inst_cellmath__220__188__I5 (.Y(N59), .A(inst_cellmath__220__188__in1[27]), .B(inst_cellmath__220__188__in1[28]), .S0(N341));
MX2XL inst_cellmath__220__188__I6 (.Y(N60), .A(inst_cellmath__220__188__in1[28]), .B(inst_cellmath__220__188__in1[29]), .S0(N341));
MX2XL inst_cellmath__220__188__I7 (.Y(N61), .A(inst_cellmath__220__188__in1[29]), .B(inst_cellmath__220__188__in1[30]), .S0(N341));
MX2XL inst_cellmath__220__188__I8 (.Y(N62), .A(inst_cellmath__220__188__in1[30]), .B(inst_cellmath__220__188__in1[31]), .S0(N341));
MX2XL inst_cellmath__220__188__I9 (.Y(N63), .A(inst_cellmath__220__188__in1[31]), .B(inst_cellmath__220__188__in1[32]), .S0(N341));
MX2XL inst_cellmath__220__188__I10 (.Y(N64), .A(inst_cellmath__220__188__in1[32]), .B(inst_cellmath__220__188__in1[33]), .S0(N341));
MX2XL inst_cellmath__220__188__I11 (.Y(N65), .A(inst_cellmath__220__188__in1[33]), .B(inst_cellmath__220__188__in1[34]), .S0(N341));
MX2XL inst_cellmath__220__188__I12 (.Y(N66), .A(inst_cellmath__220__188__in1[34]), .B(inst_cellmath__220__188__in1[35]), .S0(N341));
MX2XL inst_cellmath__220__188__I13 (.Y(N67), .A(inst_cellmath__220__188__in1[35]), .B(inst_cellmath__220__188__in1[36]), .S0(N341));
MX2XL inst_cellmath__220__188__I14 (.Y(N68), .A(inst_cellmath__220__188__in1[36]), .B(inst_cellmath__220__188__in1[37]), .S0(N341));
MX2XL inst_cellmath__220__188__I15 (.Y(N69), .A(inst_cellmath__220__188__in1[37]), .B(inst_cellmath__220__188__in1[38]), .S0(N341));
MX2XL inst_cellmath__220__188__I16 (.Y(N70), .A(inst_cellmath__220__188__in1[38]), .B(inst_cellmath__220__188__in1[39]), .S0(N341));
MX2XL inst_cellmath__220__188__I17 (.Y(N71), .A(inst_cellmath__220__188__in1[39]), .B(inst_cellmath__220__188__in1[40]), .S0(N341));
MX2XL inst_cellmath__220__188__I18 (.Y(N72), .A(inst_cellmath__220__188__in1[40]), .B(inst_cellmath__220__188__in1[41]), .S0(N341));
MX2XL inst_cellmath__220__188__I19 (.Y(N73), .A(inst_cellmath__220__188__in1[41]), .B(inst_cellmath__220__188__in1[42]), .S0(N341));
MX2XL inst_cellmath__220__188__I20 (.Y(N74), .A(inst_cellmath__220__188__in1[42]), .B(inst_cellmath__220__188__in1[43]), .S0(N341));
MX2XL inst_cellmath__220__188__I21 (.Y(N75), .A(inst_cellmath__220__188__in1[43]), .B(inst_cellmath__220__188__in1[44]), .S0(N341));
MX2XL inst_cellmath__220__188__I22 (.Y(N76), .A(inst_cellmath__220__188__in1[44]), .B(inst_cellmath__220__188__in1[45]), .S0(N341));
MX2XL inst_cellmath__220__188__I23 (.Y(N77), .A(inst_cellmath__220__188__in1[45]), .B(inst_cellmath__220__188__in1[46]), .S0(N341));
MX2XL inst_cellmath__220__188__I24 (.Y(N78), .A(inst_cellmath__220__188__in1[46]), .B(inst_cellmath__220__188__in1[47]), .S0(N341));
CLKINVX12 inst_cellmath__220__188__I258 (.Y(N342), .A(inst_cellmath__220__188__in0[1]));
NAND2XL inst_cellmath__220__188__I52 (.Y(N106), .A(N55), .B(N342));
NAND2XL inst_cellmath__220__188__I53 (.Y(N108), .A(N57), .B(N342));
MXI2XL inst_cellmath__220__188__I54 (.Y(N110), .A(N55), .B(N58), .S0(N342));
MXI2XL inst_cellmath__220__188__I55 (.Y(N111), .A(N57), .B(N59), .S0(N342));
MXI2X1 inst_cellmath__220__188__I56 (.Y(N112), .A(N58), .B(N60), .S0(N342));
MXI2X1 inst_cellmath__220__188__I57 (.Y(N113), .A(N59), .B(N61), .S0(N342));
MXI2XL inst_cellmath__220__188__I58 (.Y(N114), .A(N60), .B(N62), .S0(N342));
MXI2XL inst_cellmath__220__188__I59 (.Y(N115), .A(N61), .B(N63), .S0(N342));
MXI2XL inst_cellmath__220__188__I60 (.Y(N116), .A(N62), .B(N64), .S0(N342));
MXI2XL inst_cellmath__220__188__I61 (.Y(N117), .A(N63), .B(N65), .S0(N342));
MXI2XL inst_cellmath__220__188__I62 (.Y(N118), .A(N64), .B(N66), .S0(N342));
MXI2XL inst_cellmath__220__188__I63 (.Y(N119), .A(N65), .B(N67), .S0(N342));
MXI2XL inst_cellmath__220__188__I64 (.Y(N120), .A(N66), .B(N68), .S0(N342));
MXI2X1 inst_cellmath__220__188__I65 (.Y(N121), .A(N67), .B(N69), .S0(N342));
MXI2XL inst_cellmath__220__188__I66 (.Y(N122), .A(N68), .B(N70), .S0(N342));
MXI2XL inst_cellmath__220__188__I67 (.Y(N123), .A(N69), .B(N71), .S0(N342));
MXI2X1 inst_cellmath__220__188__I68 (.Y(N124), .A(N70), .B(N72), .S0(N342));
MXI2X1 inst_cellmath__220__188__I69 (.Y(N125), .A(N71), .B(N73), .S0(N342));
MXI2XL inst_cellmath__220__188__I70 (.Y(N126), .A(N72), .B(N74), .S0(N342));
MXI2XL inst_cellmath__220__188__I71 (.Y(N127), .A(N73), .B(N75), .S0(N342));
MXI2XL inst_cellmath__220__188__I72 (.Y(N128), .A(N74), .B(N76), .S0(N342));
MXI2XL inst_cellmath__220__188__I73 (.Y(N129), .A(N75), .B(N77), .S0(N342));
MXI2XL inst_cellmath__220__188__I74 (.Y(N130), .A(N76), .B(N78), .S0(N342));
INVX2 inst_cellmath__220__188__I259 (.Y(N343), .A(inst_cellmath__220__188__in0[2]));
INVXL inst_cellmath__220__188__I265 (.Y(N349), .A(N343));
INVX1 inst_cellmath__220__188__I264 (.Y(N348), .A(N343));
INVX2 inst_cellmath__220__188__I263 (.Y(N347), .A(N343));
NOR2XL inst_cellmath__220__188__I102 (.Y(N158), .A(N106), .B(N349));
NOR2XL inst_cellmath__220__188__I103 (.Y(N160), .A(N108), .B(N349));
NOR2XL inst_cellmath__220__188__I104 (.Y(N162), .A(N110), .B(N349));
NOR2XL inst_cellmath__220__188__I105 (.Y(N164), .A(N111), .B(N348));
MXI2X1 inst_cellmath__220__188__I106 (.Y(N166), .A(N112), .B(N106), .S0(N348));
MXI2X1 inst_cellmath__220__188__I107 (.Y(N167), .A(N113), .B(N108), .S0(N348));
MXI2XL inst_cellmath__220__188__I108 (.Y(N168), .A(N114), .B(N110), .S0(N348));
MXI2XL inst_cellmath__220__188__I109 (.Y(N169), .A(N115), .B(N111), .S0(N347));
MXI2XL inst_cellmath__220__188__I110 (.Y(N170), .A(N116), .B(N112), .S0(N347));
MXI2XL inst_cellmath__220__188__I111 (.Y(N171), .A(N117), .B(N113), .S0(N347));
MXI2XL inst_cellmath__220__188__I112 (.Y(N172), .A(N118), .B(N114), .S0(N347));
MXI2XL inst_cellmath__220__188__I113 (.Y(N173), .A(N119), .B(N115), .S0(N347));
MXI2XL inst_cellmath__220__188__I114 (.Y(N174), .A(N120), .B(N116), .S0(N347));
MXI2XL inst_cellmath__220__188__I115 (.Y(N175), .A(N121), .B(N117), .S0(N347));
MXI2XL inst_cellmath__220__188__I116 (.Y(N176), .A(N122), .B(N118), .S0(N347));
MXI2XL inst_cellmath__220__188__I117 (.Y(N177), .A(N123), .B(N119), .S0(N348));
MXI2XL inst_cellmath__220__188__I118 (.Y(N178), .A(N124), .B(N120), .S0(N348));
MXI2XL inst_cellmath__220__188__I119 (.Y(N179), .A(N125), .B(N121), .S0(N348));
MXI2XL inst_cellmath__220__188__I120 (.Y(N180), .A(N126), .B(N122), .S0(N348));
MXI2XL inst_cellmath__220__188__I121 (.Y(N181), .A(N127), .B(N123), .S0(N347));
MXI2XL inst_cellmath__220__188__I122 (.Y(N182), .A(N128), .B(N124), .S0(N347));
MXI2XL inst_cellmath__220__188__I123 (.Y(N183), .A(N129), .B(N125), .S0(N347));
MXI2XL inst_cellmath__220__188__I124 (.Y(N184), .A(N130), .B(N126), .S0(N347));
BUFX2 inst_cellmath__220__188__I283 (.Y(N351), .A(inst_cellmath__220__188__in0[4]));
INVX2 inst_cellmath__220__188__I273 (.Y(N357), .A(N351));
INVX1 inst_cellmath__220__188__I271 (.Y(N355), .A(N351));
NAND2XL inst_cellmath__220__188__I152 (.Y(N212), .A(N158), .B(N357));
NAND2XL inst_cellmath__220__188__I153 (.Y(N214), .A(N160), .B(N357));
NAND2XL inst_cellmath__220__188__I154 (.Y(N216), .A(N162), .B(N357));
NAND2XL inst_cellmath__220__188__I155 (.Y(N218), .A(N164), .B(N357));
NAND2XL inst_cellmath__220__188__I156 (.Y(N220), .A(N166), .B(N357));
NAND2XL inst_cellmath__220__188__I157 (.Y(N222), .A(N167), .B(N357));
NAND2XL inst_cellmath__220__188__I158 (.Y(N224), .A(N168), .B(N357));
NAND2XL inst_cellmath__220__188__I159 (.Y(N226), .A(N169), .B(N355));
NAND2XL inst_cellmath__220__188__I160 (.Y(N228), .A(N170), .B(N355));
NAND2XL inst_cellmath__220__188__I161 (.Y(N230), .A(N171), .B(N355));
NAND2XL inst_cellmath__220__188__I162 (.Y(N232), .A(N172), .B(N355));
NAND2XL inst_cellmath__220__188__I163 (.Y(N234), .A(N173), .B(N355));
NAND2XL inst_cellmath__220__188__I164 (.Y(N236), .A(N174), .B(N355));
NAND2XL inst_cellmath__220__188__I165 (.Y(N238), .A(N175), .B(N355));
NAND2XL inst_cellmath__220__188__I166 (.Y(N240), .A(N176), .B(N355));
NAND2XL inst_cellmath__220__188__I167 (.Y(N242), .A(N177), .B(N355));
MXI2XL inst_cellmath__220__188__I168 (.Y(N244), .A(N158), .B(N178), .S0(N355));
MXI2XL inst_cellmath__220__188__I169 (.Y(N245), .A(N160), .B(N179), .S0(N355));
MXI2XL inst_cellmath__220__188__I170 (.Y(N246), .A(N162), .B(N180), .S0(N355));
MXI2XL inst_cellmath__220__188__I171 (.Y(N247), .A(N164), .B(N181), .S0(N357));
MXI2XL inst_cellmath__220__188__I172 (.Y(N248), .A(N166), .B(N182), .S0(N357));
MXI2XL inst_cellmath__220__188__I173 (.Y(N249), .A(N167), .B(N183), .S0(N357));
MXI2XL inst_cellmath__220__188__I174 (.Y(N250), .A(N168), .B(N184), .S0(N357));
INVXL inst_cellmath__220__188__I274 (.Y(N358), .A(inst_cellmath__220__188__in0[3]));
INVX1 inst_cellmath__220__188__I280 (.Y(N364), .A(N358));
INVXL inst_cellmath__220__188__I276 (.Y(N360), .A(N358));
NOR2XL inst_cellmath__220__188__I202 (.Y(inst_cellmath__220__188__out0[0]), .A(N212), .B(N364));
NOR2XL inst_cellmath__220__188__I203 (.Y(inst_cellmath__220__188__out0[1]), .A(N214), .B(N364));
NOR2XL inst_cellmath__220__188__I204 (.Y(inst_cellmath__220__188__out0[2]), .A(N216), .B(N364));
NOR2XL inst_cellmath__220__188__I205 (.Y(inst_cellmath__220__188__out0[3]), .A(N218), .B(N364));
NOR2XL inst_cellmath__220__188__I206 (.Y(inst_cellmath__220__188__out0[4]), .A(N220), .B(N364));
NOR2XL inst_cellmath__220__188__I207 (.Y(inst_cellmath__220__188__out0[5]), .A(N222), .B(N364));
NOR2XL inst_cellmath__220__188__I208 (.Y(inst_cellmath__220__188__out0[6]), .A(N224), .B(N364));
NOR2XL inst_cellmath__220__188__I209 (.Y(inst_cellmath__220__188__out0[7]), .A(N226), .B(N364));
MXI2X1 inst_cellmath__220__188__I210 (.Y(inst_cellmath__220__188__out0[8]), .A(N228), .B(N212), .S0(N364));
MXI2X1 inst_cellmath__220__188__I211 (.Y(inst_cellmath__220__188__out0[9]), .A(N230), .B(N214), .S0(N364));
MXI2X1 inst_cellmath__220__188__I212 (.Y(inst_cellmath__220__188__out0[10]), .A(N232), .B(N216), .S0(N364));
MXI2XL inst_cellmath__220__188__I213 (.Y(inst_cellmath__220__188__out0[11]), .A(N234), .B(N218), .S0(N364));
MXI2XL inst_cellmath__220__188__I214 (.Y(inst_cellmath__220__188__out0[12]), .A(N236), .B(N220), .S0(N364));
MXI2XL inst_cellmath__220__188__I215 (.Y(inst_cellmath__220__188__out0[13]), .A(N238), .B(N222), .S0(N364));
MXI2XL inst_cellmath__220__188__I216 (.Y(inst_cellmath__220__188__out0[14]), .A(N240), .B(N224), .S0(N364));
MXI2X1 inst_cellmath__220__188__I217 (.Y(inst_cellmath__220__188__out0[15]), .A(N242), .B(N226), .S0(N360));
MXI2XL inst_cellmath__220__188__I218 (.Y(inst_cellmath__220__188__out0[16]), .A(N244), .B(N228), .S0(N360));
MXI2XL inst_cellmath__220__188__I219 (.Y(inst_cellmath__220__188__out0[17]), .A(N245), .B(N230), .S0(N360));
MXI2XL inst_cellmath__220__188__I220 (.Y(inst_cellmath__220__188__out0[18]), .A(N246), .B(N232), .S0(N360));
MXI2XL inst_cellmath__220__188__I221 (.Y(inst_cellmath__220__188__out0[19]), .A(N247), .B(N234), .S0(N360));
MXI2XL inst_cellmath__220__188__I222 (.Y(inst_cellmath__220__188__out0[20]), .A(N248), .B(N236), .S0(N360));
MXI2XL inst_cellmath__220__188__I223 (.Y(inst_cellmath__220__188__out0[21]), .A(N249), .B(N238), .S0(N360));
MXI2XL inst_cellmath__220__188__I224 (.Y(inst_cellmath__220__188__out0[22]), .A(N250), .B(N240), .S0(N360));
endmodule

module cynw_cm_float_sin_inst_cellmath__221__195__bdw1946085813_bdw (
	inst_cellmath__221__195__out0,
	inst_cellmath__221__195__in0
	); /* architecture "gate_level" */ 
output [6:0] inst_cellmath__221__195__out0;
input [4:0] inst_cellmath__221__195__in0;
INVXL inst_cellmath__221__195__I5 (.Y(inst_cellmath__221__195__out0[0]), .A(inst_cellmath__221__195__in0[0]));
INVXL inst_cellmath__221__195__I6 (.Y(inst_cellmath__221__195__out0[1]), .A(inst_cellmath__221__195__in0[1]));
INVXL inst_cellmath__221__195__I7 (.Y(inst_cellmath__221__195__out0[2]), .A(inst_cellmath__221__195__in0[2]));
INVXL inst_cellmath__221__195__I8 (.Y(inst_cellmath__221__195__out0[3]), .A(inst_cellmath__221__195__in0[3]));
INVXL inst_cellmath__221__195__I9 (.Y(inst_cellmath__221__195__out0[4]), .A(inst_cellmath__221__195__in0[4]));
assign inst_cellmath__221__195__out0[5] = 1'B1;
assign inst_cellmath__221__195__out0[6] = 1'B1;
endmodule

module cynw_cm_float_sin_inst_cellmath__220_2WWMM_bdw1946085813_bdw (
	inst_cellmath__220_2WWMM_out0,
	inst_cellmath__220_2WWMM_in0,
	inst_cellmath__220_2WWMM_in1,
	inst_cellmath__220_2WWMM_in2,
	inst_cellmath__220_2WWMM_in3,
	inst_cellmath__220_2WWMM_in4,
	inst_cellmath__220_2WWMM_in5
	); /* architecture "gate_level" */ 
output [30:0] inst_cellmath__220_2WWMM_out0;
input [6:0] inst_cellmath__220_2WWMM_in0;
input [22:0] inst_cellmath__220_2WWMM_in1;
input  inst_cellmath__220_2WWMM_in2;
input [0:0] inst_cellmath__220_2WWMM_in3;
input [22:0] inst_cellmath__220_2WWMM_in4;
input [7:0] inst_cellmath__220_2WWMM_in5;
wire N166,N168,N170,N172,N174,N176,N178 
	,N324,N410;
NOR2X1 inst_cellmath__220_2WWMM_I0 (.Y(N324), .A(inst_cellmath__220_2WWMM_in2), .B(inst_cellmath__220_2WWMM_in3[0]));
AOI22XL inst_cellmath__220_2WWMM_I6 (.Y(N166), .A0(inst_cellmath__220_2WWMM_in5[0]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[0]));
AOI22XL inst_cellmath__220_2WWMM_I7 (.Y(N168), .A0(inst_cellmath__220_2WWMM_in5[1]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[1]));
AOI22XL inst_cellmath__220_2WWMM_I8 (.Y(N170), .A0(inst_cellmath__220_2WWMM_in5[2]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[2]));
AOI22XL inst_cellmath__220_2WWMM_I9 (.Y(N172), .A0(inst_cellmath__220_2WWMM_in5[3]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[3]));
AOI22XL inst_cellmath__220_2WWMM_I10 (.Y(N174), .A0(inst_cellmath__220_2WWMM_in5[4]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[4]));
AOI22XL inst_cellmath__220_2WWMM_I11 (.Y(N176), .A0(inst_cellmath__220_2WWMM_in5[5]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[5]));
AOI22XL inst_cellmath__220_2WWMM_I12 (.Y(N178), .A0(inst_cellmath__220_2WWMM_in5[6]), .A1(inst_cellmath__220_2WWMM_in3[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in0[6]));
AND2XL inst_cellmath__220_2WWMM_I13 (.Y(inst_cellmath__220_2WWMM_out0[7]), .A(inst_cellmath__220_2WWMM_in5[7]), .B(inst_cellmath__220_2WWMM_in3[0]));
AO22XL inst_cellmath__220_2WWMM_I14 (.Y(inst_cellmath__220_2WWMM_out0[8]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[0]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[0]));
AO22XL inst_cellmath__220_2WWMM_I15 (.Y(inst_cellmath__220_2WWMM_out0[9]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[1]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[1]));
AO22XL inst_cellmath__220_2WWMM_I16 (.Y(inst_cellmath__220_2WWMM_out0[10]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[2]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[2]));
AO22XL inst_cellmath__220_2WWMM_I17 (.Y(inst_cellmath__220_2WWMM_out0[11]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[3]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[3]));
AO22XL inst_cellmath__220_2WWMM_I18 (.Y(inst_cellmath__220_2WWMM_out0[12]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[4]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[4]));
AO22XL inst_cellmath__220_2WWMM_I19 (.Y(inst_cellmath__220_2WWMM_out0[13]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[5]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[5]));
AO22XL inst_cellmath__220_2WWMM_I20 (.Y(inst_cellmath__220_2WWMM_out0[14]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[6]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[6]));
AO22XL inst_cellmath__220_2WWMM_I21 (.Y(inst_cellmath__220_2WWMM_out0[15]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[7]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[7]));
AO22XL inst_cellmath__220_2WWMM_I22 (.Y(inst_cellmath__220_2WWMM_out0[16]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[8]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[8]));
AO22XL inst_cellmath__220_2WWMM_I23 (.Y(inst_cellmath__220_2WWMM_out0[17]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[9]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[9]));
AO22XL inst_cellmath__220_2WWMM_I24 (.Y(inst_cellmath__220_2WWMM_out0[18]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[10]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[10]));
AO22XL inst_cellmath__220_2WWMM_I25 (.Y(inst_cellmath__220_2WWMM_out0[19]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[11]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[11]));
AO22XL inst_cellmath__220_2WWMM_I26 (.Y(inst_cellmath__220_2WWMM_out0[20]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[12]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[12]));
AO22XL inst_cellmath__220_2WWMM_I27 (.Y(inst_cellmath__220_2WWMM_out0[21]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[13]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[13]));
AO22XL inst_cellmath__220_2WWMM_I28 (.Y(inst_cellmath__220_2WWMM_out0[22]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[14]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[14]));
AO22XL inst_cellmath__220_2WWMM_I29 (.Y(inst_cellmath__220_2WWMM_out0[23]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[15]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[15]));
AO22XL inst_cellmath__220_2WWMM_I30 (.Y(inst_cellmath__220_2WWMM_out0[24]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[16]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[16]));
AO22XL inst_cellmath__220_2WWMM_I31 (.Y(inst_cellmath__220_2WWMM_out0[25]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[17]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[17]));
AO22XL inst_cellmath__220_2WWMM_I32 (.Y(inst_cellmath__220_2WWMM_out0[26]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[18]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[18]));
AO22XL inst_cellmath__220_2WWMM_I33 (.Y(inst_cellmath__220_2WWMM_out0[27]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[19]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[19]));
AO22XL inst_cellmath__220_2WWMM_I34 (.Y(inst_cellmath__220_2WWMM_out0[28]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[20]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[20]));
AO22XL inst_cellmath__220_2WWMM_I35 (.Y(inst_cellmath__220_2WWMM_out0[29]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[21]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[21]));
AO22XL inst_cellmath__220_2WWMM_I36 (.Y(inst_cellmath__220_2WWMM_out0[30]), .A0(inst_cellmath__220_2WWMM_in3[0]), .A1(inst_cellmath__220_2WWMM_in4[22]), .B0(N324), .B1(inst_cellmath__220_2WWMM_in1[22]));
NAND2BXL inst_cellmath__220_2WWMM_I114 (.Y(N410), .AN(inst_cellmath__220_2WWMM_in3[0]), .B(inst_cellmath__220_2WWMM_in2));
NAND2XL inst_cellmath__220_2WWMM_I71 (.Y(inst_cellmath__220_2WWMM_out0[0]), .A(N166), .B(N410));
NAND2XL inst_cellmath__220_2WWMM_I72 (.Y(inst_cellmath__220_2WWMM_out0[1]), .A(N410), .B(N168));
NAND2XL inst_cellmath__220_2WWMM_I73 (.Y(inst_cellmath__220_2WWMM_out0[2]), .A(N410), .B(N170));
NAND2XL inst_cellmath__220_2WWMM_I74 (.Y(inst_cellmath__220_2WWMM_out0[3]), .A(N410), .B(N172));
NAND2XL inst_cellmath__220_2WWMM_I75 (.Y(inst_cellmath__220_2WWMM_out0[4]), .A(N410), .B(N174));
NAND2XL inst_cellmath__220_2WWMM_I76 (.Y(inst_cellmath__220_2WWMM_out0[5]), .A(N176), .B(N410));
NAND2XL inst_cellmath__220_2WWMM_I77 (.Y(inst_cellmath__220_2WWMM_out0[6]), .A(N178), .B(N410));
endmodule

module cynw_cm_float_sin_inst_cellmath__223__208__bdw1946085813_bdw (
	inst_cellmath__223__208__out0,
	inst_cellmath__223__208__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__208__out0;
input [29:0] inst_cellmath__223__208__in0;
wire N37,N40,N42,N44,N53,N54,N55 
	,N58,N59,N61,N64,N65,N66,N67,N68 
	,N70,N72,N73,N74,N75;
OR4X1 inst_cellmath__223__208__I50 (.Y(N37), .A(inst_cellmath__223__208__in0[7]), .B(inst_cellmath__223__208__in0[5]), .C(inst_cellmath__223__208__in0[6]), .D(inst_cellmath__223__208__in0[0]));
NOR3XL inst_cellmath__223__208__I51 (.Y(N40), .A(N37), .B(inst_cellmath__223__208__in0[1]), .C(inst_cellmath__223__208__in0[2]));
NOR2XL inst_cellmath__223__208__I8 (.Y(N42), .A(inst_cellmath__223__208__in0[4]), .B(inst_cellmath__223__208__in0[3]));
NAND2XL inst_cellmath__223__208__I10 (.Y(N44), .A(N42), .B(N40));
NOR3XL inst_cellmath__223__208__I53 (.Y(N64), .A(N44), .B(inst_cellmath__223__208__in0[8]), .C(inst_cellmath__223__208__in0[15]));
NOR3XL inst_cellmath__223__208__I54 (.Y(N53), .A(inst_cellmath__223__208__in0[9]), .B(inst_cellmath__223__208__in0[10]), .C(inst_cellmath__223__208__in0[12]));
NOR2XL inst_cellmath__223__208__I21 (.Y(N54), .A(inst_cellmath__223__208__in0[23]), .B(inst_cellmath__223__208__in0[16]));
NOR2XL inst_cellmath__223__208__I22 (.Y(N55), .A(inst_cellmath__223__208__in0[17]), .B(inst_cellmath__223__208__in0[22]));
NOR3XL inst_cellmath__223__208__I55 (.Y(N68), .A(inst_cellmath__223__208__in0[13]), .B(inst_cellmath__223__208__in0[11]), .C(inst_cellmath__223__208__in0[18]));
NOR2XL inst_cellmath__223__208__I25 (.Y(N58), .A(inst_cellmath__223__208__in0[24]), .B(inst_cellmath__223__208__in0[28]));
NOR2X1 inst_cellmath__223__208__I26 (.Y(N59), .A(inst_cellmath__223__208__in0[25]), .B(inst_cellmath__223__208__in0[29]));
NOR3XL inst_cellmath__223__208__I56 (.Y(N61), .A(inst_cellmath__223__208__in0[20]), .B(inst_cellmath__223__208__in0[19]), .C(inst_cellmath__223__208__in0[27]));
OR3XL inst_cellmath__223__208__I57 (.Y(N70), .A(inst_cellmath__223__208__in0[21]), .B(inst_cellmath__223__208__in0[14]), .C(inst_cellmath__223__208__in0[26]));
NAND2XL inst_cellmath__223__208__I32 (.Y(N65), .A(N64), .B(N54));
NAND2XL inst_cellmath__223__208__I33 (.Y(N66), .A(N55), .B(N58));
NAND2XL inst_cellmath__223__208__I34 (.Y(N67), .A(N59), .B(N53));
NAND2XL inst_cellmath__223__208__I36 (.Y(N73), .A(N68), .B(N61));
NOR2XL inst_cellmath__223__208__I38 (.Y(N75), .A(N70), .B(N66));
OR2XL inst_cellmath__223__208__I39 (.Y(N72), .A(N65), .B(N67));
NOR2X1 inst_cellmath__223__208__I41 (.Y(N74), .A(N73), .B(N72));
NAND2X1 inst_cellmath__223__208__I43 (.Y(inst_cellmath__223__208__out0[0]), .A(N75), .B(N74));
endmodule

module cynw_cm_float_sin_inst_cellmath__223__207__bdw1946085813_bdw (
	inst_cellmath__223__207__out0,
	inst_cellmath__223__207__in0,
	inst_cellmath__223__207__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__207__out0;
input [24:24] inst_cellmath__223__207__in0;
input  inst_cellmath__223__207__in1;
wire N6;
INVXL inst_cellmath__223__207__I1 (.Y(N6), .A(inst_cellmath__223__207__in1));
MXI2XL inst_cellmath__223__207__I2 (.Y(inst_cellmath__223__207__out0[0]), .A(N6), .B(inst_cellmath__223__207__in1), .S0(inst_cellmath__223__207__in0[24]));
endmodule

module cynw_cm_float_sin_inst_cellmath__223__199__bdw1946085813_bdw (
	inst_cellmath__223__199__out0,
	inst_cellmath__223__199__in0,
	inst_cellmath__223__199__in1,
	inst_cellmath__223__199__in2,
	inst_cellmath__223__199__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__223__199__out0;
input  inst_cellmath__223__199__in0;
input [0:0] inst_cellmath__223__199__in1,
	inst_cellmath__223__199__in2,
	inst_cellmath__223__199__in3;
wire N7,N8,N9,N10;
NOR2XL inst_cellmath__223__199__I0 (.Y(N7), .A(inst_cellmath__223__199__in0), .B(inst_cellmath__223__199__in1[0]));
NAND2XL inst_cellmath__223__199__I1 (.Y(N8), .A(N7), .B(inst_cellmath__223__199__in3[0]));
INVXL inst_cellmath__223__199__I2 (.Y(N9), .A(N8));
NAND2X2 inst_cellmath__223__199__I3 (.Y(N10), .A(N9), .B(inst_cellmath__223__199__in2[0]));
INVX1 inst_cellmath__223__199__I4 (.Y(inst_cellmath__223__199__out0[0]), .A(N10));
endmodule

module cynw_cm_float_sin_inst_cellmath__223_0_bdw1946085813_bdw (
	inst_cellmath__223_0_out0,
	inst_cellmath__223_0_in0,
	inst_cellmath__223_0_in1,
	inst_cellmath__223_0_in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__223_0_out0;
input [0:0] inst_cellmath__223_0_in0,
	inst_cellmath__223_0_in1;
input  inst_cellmath__223_0_in2;
wire N6,N7;
INVXL inst_cellmath__223_0_I0 (.Y(N6), .A(inst_cellmath__223_0_in2));
INVXL inst_cellmath__223_0_I1 (.Y(N7), .A(inst_cellmath__223_0_in0[0]));
MXI2XL inst_cellmath__223_0_I4 (.Y(inst_cellmath__223_0_out0), .A(N7), .B(N6), .S0(inst_cellmath__223_0_in1[0]));
endmodule

module cynw_cm_float_sin_inst_cellmath__224__212__bdw1946085813_bdw (
	inst_cellmath__224__212__out0,
	inst_cellmath__224__212__in0,
	inst_cellmath__224__212__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__224__212__out0;
input  inst_cellmath__224__212__in0;
input [0:0] inst_cellmath__224__212__in1;
wire N5;
INVXL inst_cellmath__224__212__I0 (.Y(N5), .A(inst_cellmath__224__212__in0));
NAND2X2 inst_cellmath__224__212__I1 (.Y(inst_cellmath__224__212__out0[0]), .A(N5), .B(inst_cellmath__224__212__in1[0]));
endmodule

module cynw_cm_float_sin_inst_cellmath__228_0_bdw1946085813_bdw (
	inst_cellmath__228_0_out0,
	inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1,
	inst_cellmath__228_0_in2
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__228_0_out0;
input [0:0] inst_cellmath__228_0_in0,
	inst_cellmath__228_0_in1;
input [7:0] inst_cellmath__228_0_in2;
wire N81;
INVXL inst_cellmath__228_0_I23 (.Y(N81), .A(inst_cellmath__228_0_in0[0]));
AO22XL inst_cellmath__228_0_I4 (.Y(inst_cellmath__228_0_out0[0]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[0]));
AO22XL inst_cellmath__228_0_I5 (.Y(inst_cellmath__228_0_out0[1]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[1]));
AO22XL inst_cellmath__228_0_I6 (.Y(inst_cellmath__228_0_out0[2]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[2]));
AO22XL inst_cellmath__228_0_I7 (.Y(inst_cellmath__228_0_out0[3]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[3]));
AO22XL inst_cellmath__228_0_I8 (.Y(inst_cellmath__228_0_out0[4]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[4]));
AO22XL inst_cellmath__228_0_I9 (.Y(inst_cellmath__228_0_out0[5]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[5]));
AO22XL inst_cellmath__228_0_I10 (.Y(inst_cellmath__228_0_out0[6]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[6]));
AO22XL inst_cellmath__228_0_I11 (.Y(inst_cellmath__228_0_out0[7]), .A0(inst_cellmath__228_0_in0[0]), .A1(inst_cellmath__228_0_in1[0]), .B0(N81), .B1(inst_cellmath__228_0_in2[7]));
endmodule

module cynw_cm_float_sin_inst_cellmath__231_0_bdw1946085813_bdw (
	inst_cellmath__231_0_out0,
	inst_cellmath__231_0_in0,
	inst_cellmath__231_0_in1,
	inst_cellmath__231_0_in2,
	inst_cellmath__231_0_in3
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__231_0_out0;
input  inst_cellmath__231_0_in0;
input [0:0] inst_cellmath__231_0_in1;
input [30:8] inst_cellmath__231_0_in2;
input [46:46] inst_cellmath__231_0_in3;
wire N202;
INVXL inst_cellmath__231_0_I52 (.Y(N202), .A(inst_cellmath__231_0_in1[0]));
AO22XL inst_cellmath__231_0_I4 (.Y(inst_cellmath__231_0_out0[0]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[8]));
AO22XL inst_cellmath__231_0_I5 (.Y(inst_cellmath__231_0_out0[1]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[9]));
AO22XL inst_cellmath__231_0_I6 (.Y(inst_cellmath__231_0_out0[2]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[10]));
AO22XL inst_cellmath__231_0_I7 (.Y(inst_cellmath__231_0_out0[3]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[11]));
AO22XL inst_cellmath__231_0_I8 (.Y(inst_cellmath__231_0_out0[4]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[12]));
AO22XL inst_cellmath__231_0_I9 (.Y(inst_cellmath__231_0_out0[5]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[13]));
AO22XL inst_cellmath__231_0_I10 (.Y(inst_cellmath__231_0_out0[6]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[14]));
AO22XL inst_cellmath__231_0_I11 (.Y(inst_cellmath__231_0_out0[7]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[15]));
AO22XL inst_cellmath__231_0_I12 (.Y(inst_cellmath__231_0_out0[8]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[16]));
AO22XL inst_cellmath__231_0_I13 (.Y(inst_cellmath__231_0_out0[9]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[17]));
AO22XL inst_cellmath__231_0_I14 (.Y(inst_cellmath__231_0_out0[10]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[18]));
AO22XL inst_cellmath__231_0_I15 (.Y(inst_cellmath__231_0_out0[11]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[19]));
AO22XL inst_cellmath__231_0_I16 (.Y(inst_cellmath__231_0_out0[12]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[20]));
AO22XL inst_cellmath__231_0_I17 (.Y(inst_cellmath__231_0_out0[13]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[21]));
AO22XL inst_cellmath__231_0_I18 (.Y(inst_cellmath__231_0_out0[14]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[22]));
AO22XL inst_cellmath__231_0_I19 (.Y(inst_cellmath__231_0_out0[15]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[23]));
AO22XL inst_cellmath__231_0_I20 (.Y(inst_cellmath__231_0_out0[16]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[24]));
AO22XL inst_cellmath__231_0_I21 (.Y(inst_cellmath__231_0_out0[17]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[25]));
AO22XL inst_cellmath__231_0_I22 (.Y(inst_cellmath__231_0_out0[18]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[26]));
AO22XL inst_cellmath__231_0_I23 (.Y(inst_cellmath__231_0_out0[19]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[27]));
AO22XL inst_cellmath__231_0_I24 (.Y(inst_cellmath__231_0_out0[20]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[28]));
AO22XL inst_cellmath__231_0_I25 (.Y(inst_cellmath__231_0_out0[21]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[29]));
AO22XL inst_cellmath__231_0_I26 (.Y(inst_cellmath__231_0_out0[22]), .A0(inst_cellmath__231_0_in1[0]), .A1(inst_cellmath__231_0_in0), .B0(N202), .B1(inst_cellmath__231_0_in2[30]));
endmodule

/* CADENCE  vrXzTQzfqBg= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




