/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:21:38 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_cos_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__19,
	inst_cellmath__24;
wire [8:0] inst_cellmath__42;
wire [22:0] inst_cellmath__61;
wire  inst_cellmath__68;
wire [0:0] inst_cellmath__115__W1;
wire [29:0] inst_cellmath__195;
wire [20:0] inst_cellmath__197;
wire [32:0] inst_cellmath__198;
wire [49:0] inst_cellmath__201;
wire [46:0] inst_cellmath__203__W0, inst_cellmath__203__W1;
wire [30:0] inst_cellmath__210;
wire [4:0] inst_cellmath__215;
wire N493,N548,N549,N550,N551,N585,N594 
	,N595,N623,N624,N625,N626,N627,N628,N630 
	,N631,N632,N633,N634,N635,N636,N637,N638 
	,N639,N640,N641,N642,N643,N644,N645,N646 
	,N647,N648,N649,N650,N651,N652,N665,N666 
	,N667,N668,N669,N670,N671,N672,N673,N674 
	,N675,N677,N678,N679,N680,N681,N682,N683 
	,N684,N685,N686,N687,N688,N689,N690,N691 
	,N692,N693,N694,N696,N697,N698,N699,N700 
	,N701,N702,N703,N704,N705,N706,N707,N708 
	,N709,N710,N711,N712,N713,N741,N753,N761 
	,N3808,N3809,N3810,N5559,N5560,N5561,N5562,N5563 
	,N5564,N5565,N5566,N5569,N5570,N5572,N5573,N5574 
	,N5575,N5576,N5577,N5578,N5580,N5581,N5582,N5583 
	,N5587,N5588,N5589,N5590,N5591,N5592,N5594,N5595 
	,N5597,N5598,N5600,N5601,N5602,N5603,N5604,N5605 
	,N5606,N5607,N5608,N5609,N5610,N5611,N5614,N5615 
	,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623 
	,N5624,N5626,N5627,N5628,N5629,N5630,N5631,N5634 
	,N5635,N5637,N5638,N5639,N5640,N5641,N5643,N5644 
	,N5645,N5646,N5647,N5648,N5649,N5650,N5651,N5652 
	,N5653,N5655,N5656,N5657,N5658,N5659,N5660,N5662 
	,N5663,N5664,N5666,N5668,N5669,N5671,N5672,N5673 
	,N5674,N5675,N5677,N5678,N5679,N5680,N5681,N5682 
	,N5683,N5685,N5686,N5687,N5688,N5689,N5691,N5693 
	,N5694,N5695,N5698,N5699,N5700,N5701,N5702,N5703 
	,N5704,N5705,N5706,N5707,N5708,N5710,N5711,N5712 
	,N5713,N5716,N5717,N5718,N5720,N5721,N5723,N5725 
	,N5726,N5727,N5729,N5730,N5731,N5732,N5733,N5734 
	,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742 
	,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751 
	,N5752,N5753,N5754,N5755,N5757,N5758,N5759,N5763 
	,N5766,N5767,N5768,N5769,N5770,N5771,N5772,N5773 
	,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781 
	,N5784,N5785,N5786,N5787,N5788,N5789,N5792,N5793 
	,N5795,N5798,N5799,N5801,N5802,N5803,N5804,N5806 
	,N5808,N5809,N5810,N5813,N5814,N5815,N5816,N5817 
	,N5818,N5819,N5820,N5821,N5823,N5824,N5825,N5827 
	,N5828,N5829,N5830,N5832,N5833,N5834,N5835,N5836 
	,N5837,N5838,N5839,N5840,N5842,N5843,N5844,N5846 
	,N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854 
	,N5855,N5856,N5857,N5861,N5862,N5865,N5866,N5867 
	,N5868,N5869,N5870,N5871,N5872,N5875,N5876,N5878 
	,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5889 
	,N5890,N5891,N5893,N5894,N5895,N5896,N5897,N5898 
	,N5899,N5901,N5902,N5903,N5905,N5906,N5909,N5910 
	,N5911,N5912,N5914,N5915,N5916,N5917,N5918,N5919 
	,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928 
	,N5929,N5932,N5933,N5934,N5935,N5936,N5937,N5940 
	,N5941,N5942,N5944,N5945,N5946,N5947,N5949,N5950 
	,N5952,N5954,N5955,N5956,N5957,N5958,N5959,N5960 
	,N5961,N5962,N5965,N5966,N5968,N5969,N5970,N5971 
	,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980 
	,N5981,N5982,N5983,N5984,N5987,N5988,N5989,N5991 
	,N5993,N5995,N5997,N5998,N6001,N6002,N6003,N6004 
	,N6005,N6006,N6007,N6009,N6010,N6012,N6013,N6014 
	,N6015,N6017,N6018,N6019,N6020,N6021,N6022,N6023 
	,N6025,N6026,N6029,N6030,N6032,N6033,N6034,N6035 
	,N6036,N6037,N6038,N6040,N6041,N6044,N6045,N6046 
	,N6048,N6049,N6050,N6051,N6052,N6053,N6054,N6055 
	,N6056,N6058,N6060,N6063,N6064,N6065,N6068,N6069 
	,N6070,N6071,N6072,N6073,N6075,N6077,N6078,N6079 
	,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089 
	,N6090,N6091,N6092,N6094,N6095,N6096,N6097,N6099 
	,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107 
	,N6108,N6109,N6110,N6111,N6112,N6114,N6115,N6116 
	,N6117,N6118,N6119,N6120,N6122,N6123,N6124,N6126 
	,N6127,N6130,N6131,N6132,N6133,N6134,N6135,N6136 
	,N6137,N6138,N6140,N6141,N6142,N6143,N6144,N6146 
	,N6147,N6148,N6150,N6151,N6152,N6153,N6154,N6155 
	,N6156,N6157,N6158,N6162,N6163,N6164,N6166,N6167 
	,N6168,N6169,N6170,N6171,N6172,N6173,N6174,N6175 
	,N6176,N6179,N6180,N6181,N6182,N6183,N6184,N6186 
	,N6188,N6189,N6190,N6191,N6192,N6194,N6195,N6196 
	,N6197,N6198,N6199,N6200,N6201,N6203,N6204,N6206 
	,N6207,N6208,N6210,N6211,N6212,N6213,N6214,N6215 
	,N6216,N6217,N6218,N6219,N6220,N6222,N6223,N6224 
	,N6225,N6226,N6227,N6228,N6230,N6232,N6233,N6234 
	,N6235,N6236,N6237,N6239,N6240,N6241,N6242,N6243 
	,N6244,N6245,N6246,N6247,N6248,N6250,N6251,N6254 
	,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6263 
	,N6265,N6266,N6267,N6270,N6271,N6272,N6274,N6275 
	,N6276,N6277,N6278,N6279,N6281,N6283,N6284,N6285 
	,N6286,N6288,N6289,N6290,N6291,N6292,N6296,N6297 
	,N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306 
	,N6307,N6308,N6309,N6310,N6311,N6313,N6314,N6315 
	,N6317,N6318,N6319,N6320,N6321,N6322,N6325,N6326 
	,N6327,N6330,N6333,N6334,N6335,N6336,N6337,N6338 
	,N6339,N6341,N6342,N6343,N6345,N6346,N6347,N6348 
	,N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356 
	,N6357,N6358,N6359,N6363,N6366,N6368,N6369,N6370 
	,N6371,N6373,N6374,N6376,N6377,N6378,N6379,N6380 
	,N6381,N6382,N6385,N6386,N6387,N6388,N6389,N6390 
	,N6391,N6392,N6393,N6394,N6395,N6396,N6398,N6399 
	,N6400,N6401,N6403,N6404,N6405,N6406,N6407,N6408 
	,N6409,N6410,N6412,N6413,N6414,N6415,N6416,N6418 
	,N6419,N6420,N6421,N7264,N7267,N7268,N7270,N7271 
	,N7280,N7281,N7284,N7287,N7289,N7291,N7293,N7318 
	,N7320,N7321,N7322,N7324,N7325,N7329,N7331,N7332 
	,N7333,N7335,N7337,N7341,N7343,N7344,N7346,N7348 
	,N7349,N7351,N7353,N7354,N7355,N7357,N7360,N7362 
	,N7363,N7365,N7366,N7368,N7370,N7372,N7373,N7375 
	,N7376,N7378,N7379,N7381,N7385,N7387,N7388,N7390 
	,N7391,N7392,N7394,N7395,N7398,N7400,N7401,N7402 
	,N7404,N7407,N7408,N7410,N7411,N7412,N7414,N7416 
	,N7418,N7419,N7421,N7423,N7424,N7426,N7428,N7431 
	,N7432,N7434,N7436,N7437,N7438,N7441,N7443,N7444 
	,N7446,N7447,N7448,N7450,N7453,N7454,N7456,N7457 
	,N7460,N7462,N7463,N7464,N7466,N7467,N7468,N7469 
	,N7472,N7473,N7475,N7477,N7478,N7480,N7484,N7486 
	,N7487,N7489,N7492,N7494,N7495,N7496,N7498,N7499 
	,N7501,N7503,N7506,N7507,N7508,N7510,N7512,N7513 
	,N7516,N7518,N7519,N7521,N7522,N7524,N7525,N7528 
	,N7529,N7531,N7532,N7533,N7535,N7536,N7541,N7543 
	,N7544,N7546,N7547,N7549,N7551,N7552,N7554,N7555 
	,N7557,N7559,N7562,N7563,N7565,N7566,N7568,N7570 
	,N7809,N7812,N7833,N7882,N7883,N7884,N7885,N7886 
	,N7887,N7888,N7890,N7892,N7893,N7895,N7896,N7897 
	,N7898,N7899,N7901,N7902,N7903,N7905,N7906,N7907 
	,N7908,N7909,N7910,N7911,N7912,N7913,N7914,N7915 
	,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925 
	,N7926,N7927,N7929,N7930,N7932,N7933,N7934,N7937 
	,N7938,N7940,N7941,N7943,N7945,N7946,N7947,N7948 
	,N7949,N7950,N7951,N7952,N7953,N7957,N7958,N7959 
	,N7960,N7961,N7962,N7963,N7965,N7966,N7967,N7968 
	,N7970,N7971,N7973,N7974,N7976,N7977,N7978,N7980 
	,N7981,N7983,N7984,N7985,N7986,N7988,N7989,N7990 
	,N7991,N7993,N7994,N7995,N7996,N7997,N7998,N7999 
	,N8000,N8001,N8002,N8003,N8005,N8006,N8007,N8008 
	,N8009,N8010,N8011,N8012,N8013,N8014,N8016,N8017 
	,N8018,N8021,N8022,N8023,N8024,N8026,N8028,N8029 
	,N8030,N8031,N8033,N8034,N8035,N8037,N8038,N8039 
	,N8040,N8042,N8043,N8044,N8045,N8046,N8048,N8049 
	,N8050,N8051,N8052,N8053,N8055,N8056,N8057,N8058 
	,N8060,N8061,N8063,N8064,N8065,N8066,N8067,N8070 
	,N8071,N8073,N8074,N8075,N8076,N8077,N8079,N8080 
	,N8081,N8082,N8083,N8084,N8085,N8086,N8089,N8090 
	,N8091,N8094,N8095,N8096,N8097,N8098,N8099,N8101 
	,N8102,N8103,N8104,N8106,N8107,N8108,N8109,N8110 
	,N8112,N8113,N8114,N8116,N8117,N8120,N8121,N8122 
	,N8123,N8124,N8125,N8126,N8127,N8128,N8130,N8132 
	,N8133,N8135,N8136,N8137,N8138,N8142,N8144,N8146 
	,N8147,N8148,N8150,N8151,N8153,N8154,N8155,N8157 
	,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165 
	,N8166,N8167,N8169,N8170,N8171,N8172,N8173,N8174 
	,N8175,N8176,N8178,N8179,N8180,N8181,N8182,N8183 
	,N8184,N8185,N8186,N8187,N8188,N8191,N8192,N8194 
	,N8195,N8196,N8197,N8199,N8200,N8201,N8202,N8203 
	,N8204,N8205,N8206,N8207,N8208,N8209,N8210,N8212 
	,N8213,N8214,N8215,N8216,N8218,N8219,N8220,N8221 
	,N8222,N8223,N8227,N8231,N8232,N8233,N8234,N8236 
	,N8237,N8238,N8241,N8242,N8243,N8244,N8245,N8247 
	,N8248,N8250,N8251,N8252,N8254,N8259,N8260,N8261 
	,N8262,N8263,N8264,N8266,N8267,N8268,N8269,N8270 
	,N8271,N8272,N8273,N8274,N8275,N8276,N8277,N8279 
	,N8280,N8281,N8282,N8283,N8286,N8287,N8288,N8289 
	,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297 
	,N8300,N8302,N8303,N8304,N8305,N8306,N8307,N8308 
	,N8309,N8312,N8313,N8315,N8316,N8317,N8318,N8319 
	,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327 
	,N8328,N8329,N8330,N8331,N8333,N8334,N8335,N8336 
	,N8338,N8340,N8342,N8343,N8344,N8345,N8346,N8348 
	,N8349,N8350,N8351,N8352,N8353,N8355,N8357,N8360 
	,N8361,N8362,N8363,N8364,N8365,N8368,N8369,N8370 
	,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378 
	,N8379,N8380,N8382,N8383,N8384,N8386,N8388,N8389 
	,N8390,N8392,N8393,N8394,N8395,N8396,N8397,N8398 
	,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8407 
	,N8408,N8409,N8410,N8411,N8413,N8414,N8415,N8416 
	,N8418,N8419,N8420,N8421,N8422,N8423,N8425,N8426 
	,N8427,N8428,N8429,N8432,N8433,N8434,N8435,N8436 
	,N8437,N8439,N8440,N8441,N8442,N8444,N8445,N8446 
	,N8448,N8451,N8452,N8453,N8454,N8455,N8456,N8457 
	,N8458,N8459,N8460,N8461,N8462,N8463,N8464,N8465 
	,N8467,N8468,N8469,N8471,N8472,N8473,N8474,N8477 
	,N8478,N8479,N8480,N8481,N8483,N8484,N8485,N8488 
	,N8489,N8491,N8492,N8494,N8495,N8496,N8497,N8498 
	,N8499,N8501,N8502,N8503,N8504,N8505,N8506,N8507 
	,N8508,N8511,N8512,N8513,N8514,N8515,N8516,N8517 
	,N8519,N8520,N8522,N8523,N8524,N8525,N8526,N8527 
	,N8528,N8530,N8531,N8532,N8533,N8534,N8535,N8536 
	,N8537,N8538,N8539,N8540,N8543,N8544,N8545,N8548 
	,N8549,N8550,N8551,N8552,N8553,N8554,N8555,N8560 
	,N8562,N8563,N8564,N8565,N8566,N8568,N8569,N8571 
	,N8572,N8574,N8575,N8576,N8579,N8580,N8582,N8583 
	,N8584,N8586,N8587,N8588,N8589,N8590,N8592,N8593 
	,N8594,N8595,N8596,N8597,N8598,N8603,N8604,N8605 
	,N8606,N8607,N8608,N8609,N8610,N8611,N8612,N8613 
	,N8614,N8615,N8616,N8618,N8619,N8620,N8621,N8622 
	,N8624,N8625,N8626,N8627,N8628,N8630,N8631,N8632 
	,N8633,N8634,N8635,N8636,N8638,N8639,N8640,N8643 
	,N8644,N8645,N8646,N8647,N8648,N8650,N8651,N8652 
	,N8653,N8654,N8655,N8656,N8657,N8658,N8659,N8660 
	,N8662,N8663,N8665,N8666,N8668,N8669,N8670,N8671 
	,N8672,N8673,N8674,N8675,N8676,N8677,N8678,N8679 
	,N8680,N8682,N8683,N8684,N8685,N8686,N8687,N8689 
	,N8692,N8693,N8694,N8695,N8696,N8697,N8699,N8700 
	,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708 
	,N8709,N8711,N8712,N8713,N8714,N8715,N8717,N8719 
	,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727 
	,N8728,N8730,N8732,N8733,N8734,N8735,N8736,N8739 
	,N8741,N8743,N8744,N8745,N8747,N8748,N8749,N8750 
	,N8751,N8752,N8753,N8755,N8756,N8758,N8759,N8761 
	,N8762,N8763,N8764,N8766,N8767,N8770,N8771,N8772 
	,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780 
	,N8781,N8782,N8783,N8784,N8785,N8786,N8788,N8789 
	,N8790,N8793,N8794,N8795,N8796,N8798,N8799,N8800 
	,N8801,N8802,N8803,N8804,N8805,N8806,N8808,N8809 
	,N8811,N8812,N8813,N8815,N8816,N8817,N8819,N8820 
	,N8821,N8823,N8824,N8825,N8826,N8827,N8828,N8829 
	,N8831,N8832,N8834,N8835,N8837,N8838,N8839,N8841 
	,N8842,N8843,N8844,N8845,N8846,N8847,N8848,N8849 
	,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858 
	,N8859,N8860,N8862,N8864,N8865,N8867,N8868,N8870 
	,N8872,N8873,N8874,N8875,N8876,N8877,N8879,N8880 
	,N8881,N8884,N8886,N8887,N8888,N8890,N8891,N8892 
	,N8893,N8895,N8896,N8897,N8898,N8899,N8900,N8901 
	,N8903,N8904,N8905,N8906,N8907,N8908,N8909,N8911 
	,N8912,N8913,N8914,N8916,N8917,N8919,N8920,N8921 
	,N8922,N8923,N8924,N8925,N8927,N8928,N8930,N8931 
	,N8932,N8933,N8934,N8935,N8936,N8938,N8939,N8940 
	,N8941,N8943,N8944,N8946,N8947,N8948,N8949,N8950 
	,N8951,N8952,N8953,N8955,N8956,N8957,N8958,N8960 
	,N8962,N8963,N8964,N8966,N8967,N8968,N8969,N8970 
	,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978 
	,N8980,N8981,N8982,N8983,N8985,N8986,N8987,N8990 
	,N8991,N8992,N8994,N8995,N8997,N8998,N8999,N9002 
	,N9003,N9004,N9005,N9007,N9008,N9009,N9010,N9012 
	,N9013,N9014,N9015,N9017,N9019,N9020,N9022,N9023 
	,N9024,N9025,N9026,N9027,N9028,N9029,N9030,N9032 
	,N9033,N9034,N9035,N9036,N9037,N9041,N9042,N9043 
	,N9044,N9045,N9046,N9048,N9050,N9051,N9052,N9053 
	,N9055,N9056,N9059,N9060,N9061,N9062,N9063,N9064 
	,N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9073 
	,N9074,N9075,N9076,N9077,N9079,N9080,N9081,N9084 
	,N9085,N9086,N9087,N9089,N9090,N9091,N9092,N9093 
	,N9095,N9096,N9097,N9098,N9099,N9101,N9102,N9103 
	,N9104,N9105,N9106,N9109,N9110,N9111,N9113,N9115 
	,N9116,N9117,N9119,N9121,N9122,N9123,N9124,N9125 
	,N9126,N9127,N9128,N9130,N9131,N9132,N9133,N9134 
	,N9135,N9138,N9139,N9140,N9141,N9142,N10398,N10399 
	,N10400,N10401,N10402,N10403,N10406,N10407,N10408,N10410 
	,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418 
	,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428 
	,N10430,N10431,N10432,N10433,N10434,N10435,N10436,N10438 
	,N10439,N10440,N10441,N10442,N10443,N10444,N10445,N10447 
	,N10449,N10450,N10451,N10452,N10453,N10454,N10455,N10457 
	,N10458,N10459,N10460,N10461,N10462,N10463,N10464,N10465 
	,N10467,N10468,N10469,N10470,N10471,N10472,N10475,N10476 
	,N10477,N10478,N10479,N10480,N10481,N10483,N10484,N10486 
	,N10487,N10489,N10490,N10491,N10492,N10493,N10495,N10496 
	,N10497,N10498,N10499,N10500,N10502,N10504,N10505,N10509 
	,N10510,N10511,N10512,N10513,N10514,N10515,N10516,N10517 
	,N10518,N10519,N10520,N10523,N10525,N10527,N10528,N10529 
	,N10530,N10533,N10534,N10536,N10538,N10539,N10540,N10541 
	,N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549 
	,N10550,N10551,N10552,N10554,N10556,N10557,N10558,N10560 
	,N10561,N10562,N10565,N10566,N10568,N10569,N10572,N10573 
	,N10574,N10575,N10576,N10577,N10579,N10581,N10582,N10583 
	,N10584,N10585,N10586,N10587,N10588,N10590,N10591,N10592 
	,N10593,N10595,N10596,N10597,N10598,N10599,N10600,N10601 
	,N10603,N10604,N10605,N10606,N10608,N10609,N10610,N10611 
	,N10613,N10616,N10617,N10618,N10619,N10620,N10621,N10622 
	,N10623,N10625,N10626,N10627,N10628,N10629,N10630,N10631 
	,N10633,N10634,N10635,N10636,N10637,N10638,N10639,N10640 
	,N10644,N10645,N10648,N10649,N10650,N10651,N10652,N10653 
	,N10654,N10655,N10656,N10658,N10659,N10660,N10661,N10663 
	,N10665,N10666,N10667,N10670,N10671,N10672,N10673,N10674 
	,N10675,N10676,N10678,N10679,N10680,N10681,N10682,N10683 
	,N10684,N10686,N10687,N10688,N10690,N10691,N10692,N10693 
	,N10694,N10697,N10698,N10699,N10700,N10701,N10702,N10703 
	,N10704,N10705,N10706,N10708,N10709,N10710,N10711,N10712 
	,N10713,N10714,N10715,N10716,N10717,N10718,N10720,N10721 
	,N10722,N10723,N10724,N10725,N10726,N10727,N10728,N10729 
	,N10731,N10732,N10733,N10734,N10736,N10737,N10739,N10740 
	,N10743,N10745,N10746,N10747,N10748,N10749,N10750,N10753 
	,N10754,N10755,N10756,N10757,N10758,N10759,N10760,N10761 
	,N10763,N10764,N10765,N10768,N10773,N10774,N10775,N10776 
	,N10777,N10778,N10780,N10781,N10782,N10784,N10785,N10786 
	,N10787,N10788,N10789,N10790,N10791,N10792,N10793,N10794 
	,N10796,N10797,N10798,N10800,N10801,N10802,N10803,N10804 
	,N10805,N10807,N10808,N10809,N10810,N10811,N10812,N10813 
	,N10814,N10815,N10816,N10817,N10818,N10819,N10820,N10822 
	,N10823,N10824,N10825,N10827,N10828,N10829,N10832,N10833 
	,N10836,N10837,N10838,N10839,N10840,N10841,N10842,N10843 
	,N10845,N10847,N10848,N10849,N10850,N10851,N10852,N10853 
	,N10854,N10855,N10857,N10858,N10859,N10860,N10861,N10862 
	,N10863,N10864,N10865,N10867,N10870,N10871,N10872,N10873 
	,N10874,N10875,N10876,N10877,N10878,N10879,N10880,N10881 
	,N10882,N10883,N10885,N10887,N10888,N10889,N10890,N10891 
	,N10892,N10893,N10894,N10895,N10897,N10898,N10899,N10900 
	,N10902,N10903,N10906,N10907,N10908,N10909,N10911,N10913 
	,N10916,N10917,N10918,N10920,N10921,N10922,N10923,N10925 
	,N10926,N10927,N10928,N10930,N10932,N10933,N10935,N10936 
	,N10937,N10939,N10940,N10941,N10942,N10943,N10944,N10945 
	,N10946,N10947,N10949,N10950,N10951,N10952,N10953,N10954 
	,N10955,N10957,N10958,N10960,N10961,N10962,N10966,N10967 
	,N10968,N10969,N10970,N10971,N10972,N10973,N10974,N10975 
	,N10978,N10979,N10980,N10981,N10982,N10984,N10986,N10987 
	,N10988,N10990,N10991,N10992,N10994,N10995,N10996,N11000 
	,N11001,N11004,N11005,N11006,N11007,N11008,N11009,N11010 
	,N11011,N11013,N11014,N11015,N11016,N11017,N11018,N11019 
	,N11020,N11021,N11022,N11023,N11024,N11026,N11027,N11028 
	,N11029,N11033,N11034,N11035,N11036,N11037,N11038,N11667 
	,N11668,N11669,N11670,N11671,N11672,N11673,N11675,N11676 
	,N11677,N11679,N11680,N11681,N11682,N11683,N11684,N11685 
	,N11686,N11687,N11688,N11689,N11690,N11691,N11692,N11693 
	,N11694,N11695,N11696,N11697,N11699,N11700,N11701,N11702 
	,N11703,N11704,N11705,N11706,N11707,N11708,N11710,N11711 
	,N11712,N11715,N11716,N11717,N11718,N11719,N11720,N11721 
	,N11722,N11723,N11724,N11725,N11727,N11728,N11729,N11730 
	,N11731,N11732,N11734,N11735,N11737,N11738,N11739,N11740 
	,N11741,N11742,N11743,N11744,N11745,N11746,N11747,N11749 
	,N11750,N11751,N11752,N11753,N11755,N11756,N11757,N11758 
	,N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766 
	,N11767,N11768,N11769,N11770,N11771,N11772,N11773,N11774 
	,N11775,N11776,N11778,N11779,N11781,N11782,N11783,N11784 
	,N11785,N11786,N11787,N11788,N11790,N11791,N11792,N11793 
	,N11794,N11795,N11796,N11799,N11800,N11801,N11802,N11803 
	,N11804,N11805,N11806,N11807,N11808,N11809,N11810,N11811 
	,N11812,N11813,N11814,N11815,N11817,N11818,N11819,N11820 
	,N11821,N11822,N11823,N11824,N11826,N11827,N11828,N11829 
	,N11830,N11831,N11832,N11833,N11834,N11835,N11836,N11837 
	,N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846 
	,N11847,N11848,N11849,N11851,N11852,N11853,N11854,N11855 
	,N11856,N11857,N11858,N11859,N11862,N11863,N11864,N11865 
	,N11866,N11867,N11869,N11870,N11871,N11872,N11873,N11874 
	,N11875,N11876,N11877,N11879,N11880,N11881,N11882,N11883 
	,N11884,N11885,N11887,N11888,N11890,N11891,N11892,N11893 
	,N11894,N11895,N11896,N11897,N11898,N11899,N11901,N11902 
	,N11903,N11904,N11905,N11906,N11907,N11908,N11909,N11910 
	,N11911,N11912,N11913,N11914,N11915,N11916,N11918,N11919 
	,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927 
	,N11929,N11930,N11931,N11932,N11933,N11934,N11936,N11937 
	,N11938,N11939,N11940,N11941,N11942,N11943,N11944,N11946 
	,N11947,N11948,N11950,N11951,N11952,N11953,N11954,N11956 
	,N11957,N11959,N11960,N11961,N11962,N11963,N11964,N11965 
	,N11966,N11967,N11968,N11969,N11970,N11971,N11972,N11973 
	,N11974,N11976,N11978,N11979,N11980,N11981,N11983,N11985 
	,N11986,N11987,N11988,N11989,N11990,N11991,N11992,N11993 
	,N11994,N11995,N11996,N11997,N11998,N11999,N12000,N12002 
	,N12003,N12004,N12005,N12006,N12007,N12008,N12009,N12010 
	,N12011,N12013,N12014,N12015,N12016,N12017,N12021,N12022 
	,N12023,N12024,N12025,N12026,N12027,N12028,N12029,N12030 
	,N12031,N12032,N12033,N12034,N12035,N12036,N12037,N12038 
	,N12039,N12040,N12041,N12042,N12044,N12045,N12046,N12047 
	,N12048,N12049,N12051,N12052,N12053,N12054,N12056,N12057 
	,N12058,N12059,N12060,N12061,N12062,N12063,N12064,N12065 
	,N12066,N12067,N12068,N12069,N12070,N12071,N12072,N12073 
	,N12074,N12075,N12077,N12078,N12079,N12080,N12081,N12082 
	,N12083,N12084,N12086,N12087,N12088,N12089,N12091,N12092 
	,N12093,N12094,N12095,N12096,N12097,N12098,N12099,N12100 
	,N12101,N12103,N12104,N12105,N12106,N12108,N12109,N12110 
	,N12112,N12113,N12114,N12115,N12116,N12117,N12118,N12119 
	,N12120,N12121,N12122,N12123,N12124,N12125,N12126,N12127 
	,N12128,N12129,N12130,N12131,N12133,N12134,N12135,N12136 
	,N12137,N12138,N12139,N12140,N12141,N12142,N12143,N12144 
	,N12145,N12146,N12147,N12148,N12150,N12151,N12152,N12153 
	,N12154,N12155,N12156,N12157,N12159,N12160,N12161,N12162 
	,N12164,N12165,N12166,N12167,N12169,N12170,N12171,N12172 
	,N12173,N12174,N12175,N12176,N12177,N12178,N12179,N12180 
	,N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188 
	,N12189,N12190,N12192,N12193,N12194,N12195,N12196,N12198 
	,N12199,N12200,N12201,N12202,N12203,N12204,N12205,N12206 
	,N12207,N12208,N12209,N12211,N12212,N12213,N12214,N12215 
	,N12216,N12217,N12218,N12219,N12220,N12221,N12223,N12224 
	,N12225,N12226,N12227,N12229,N12231,N12232,N12233,N12234 
	,N12235,N12236,N12237,N12238,N12239,N12240,N12241,N12242 
	,N12243,N12244,N12245,N12246,N12247,N12248,N12249,N12250 
	,N12251,N12253,N12254,N12255,N12256,N12259,N12261,N12262 
	,N12263,N12264,N12265,N12266,N12267,N12269,N12270,N12271 
	,N12272,N12273,N12274,N12275,N12276,N12277,N12279,N12280 
	,N12281,N12282,N12283,N12284,N12285,N12287,N12288,N12289 
	,N12290,N12291,N12292,N12294,N12295,N12296,N12297,N12298 
	,N12299,N12303,N12304,N12305,N12306,N12307,N12308,N12309 
	,N12310,N12311,N12312,N12313,N12314,N12316,N12317,N12318 
	,N12319,N12321,N12323,N12324,N12325,N12326,N12327,N12328 
	,N12329,N12330,N12331,N12332,N12333,N12334,N12335,N12336 
	,N12337,N12338,N12339,N12340,N12342,N12343,N12344,N12347 
	,N12348,N12349,N12350,N12351,N12352,N12353,N12354,N12355 
	,N12356,N12357,N12358,N12359,N12361,N12362,N12363,N12364 
	,N12365,N12366,N12367,N12368,N12369,N12370,N12371,N12372 
	,N12373,N12374,N12375,N12377,N12378,N12380,N12381,N12384 
	,N12385,N12386,N12387,N12388,N12389,N12390,N12391,N12392 
	,N12393,N12394,N12395,N12396,N12397,N12398,N12399,N12400 
	,N12401,N12404,N12405,N12406,N12407,N12409,N12410,N12411 
	,N12412,N12414,N12415,N12416,N12417,N12418,N12419,N12420 
	,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428 
	,N12429,N12430,N12431,N12432,N12433,N12434,N12435,N12437 
	,N12438,N12439,N12440,N12441,N12443,N12444,N12447,N12448 
	,N12449,N12450,N12451,N12452,N12453,N12454,N12455,N12456 
	,N12457,N12458,N12459,N12460,N12461,N12462,N12463,N12464 
	,N12465,N12467,N12468,N12469,N12470,N12472,N12474,N12475 
	,N12476,N12477,N12478,N12479,N12480,N12481,N12482,N12483 
	,N12484,N12485,N12486,N12487,N12488,N12489,N12490,N12491 
	,N12492,N12493,N12495,N12496,N12497,N12498,N12499,N12501 
	,N12502,N12503,N12504,N12505,N12506,N12507,N12509,N12510 
	,N12511,N12512,N12514,N12515,N12516,N12517,N12518,N12519 
	,N12520,N12521,N12522,N12523,N12524,N12525,N12526,N12527 
	,N12528,N12529,N12531,N12532,N12533,N12534,N12536,N12537 
	,N12538,N12540,N12541,N12542,N12543,N12544,N12545,N12546 
	,N12547,N12548,N12549,N12550,N12551,N12552,N12553,N12554 
	,N12555,N12556,N12557,N12559,N12560,N12561,N12562,N12563 
	,N12564,N12566,N12567,N12568,N12569,N12570,N12571,N12572 
	,N12573,N12574,N12575,N12577,N12578,N12579,N12580,N12581 
	,N12582,N12583,N12584,N12585,N12586,N12587,N12588,N12589 
	,N12590,N12591,N12592,N12593,N12595,N12596,N12599,N12600 
	,N12601,N12602,N12603,N12604,N12605,N12606,N12607,N12608 
	,N12609,N12610,N12611,N12612,N12613,N12614,N12615,N12617 
	,N12618,N12619,N12620,N12622,N12625,N12626,N12627,N12628 
	,N12629,N12630,N12632,N12633,N12635,N12636,N12637,N12638 
	,N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646 
	,N12647,N12648,N12649,N12651,N12652,N12653,N12654,N12655 
	,N12656,N12658,N12659,N12660,N12661,N12664,N12665,N12666 
	,N12667,N12668,N12669,N12670,N12671,N12673,N12675,N12676 
	,N12677,N12679,N12680,N12682,N12683,N12684,N12685,N12686 
	,N12687,N12688,N12689,N12690,N12691,N12692,N12693,N12694 
	,N12695,N12696,N12697,N12698,N12700,N12702,N12703,N12704 
	,N12705,N12706,N12707,N12708,N12709,N12710,N12711,N12712 
	,N12713,N12714,N12716,N12717,N12718,N12719,N12720,N12721 
	,N12722,N12723,N12724,N12725,N12726,N12727,N12729,N12730 
	,N12732,N12734,N12736,N12737,N12738,N12739,N12740,N12741 
	,N12742,N12743,N12744,N12745,N12746,N12747,N12748,N12749 
	,N12750,N12751,N12752,N12755,N12756,N12757,N12758,N12759 
	,N12761,N12762,N12763,N12764,N12765,N12766,N12767,N12768 
	,N12769,N12770,N12771,N12772,N12773,N12774,N12775,N12776 
	,N12777,N12778,N12779,N12780,N12781,N12783,N12784,N12785 
	,N12786,N12787,N12789,N12791,N12792,N12793,N12794,N12795 
	,N12796,N12797,N12798,N12799,N12800,N12801,N12802,N12803 
	,N12804,N12805,N12807,N12808,N12809,N12810,N12811,N12812 
	,N12814,N12816,N12817,N12818,N12819,N12820,N12821,N12822 
	,N12823,N12824,N12825,N12826,N12827,N12828,N12829,N12830 
	,N12832,N12833,N12834,N12835,N12836,N12837,N12838,N12840 
	,N12841,N12842,N12843,N12844,N12845,N12846,N12848,N12849 
	,N12850,N12852,N12853,N12854,N12855,N12856,N12857,N12858 
	,N12859,N12860,N12861,N12862,N12863,N12864,N12866,N12867 
	,N12868,N12869,N12870,N12871,N12873,N12874,N12875,N12876 
	,N12877,N12879,N12880,N12881,N12882,N12883,N12884,N12885 
	,N12886,N12888,N12889,N12891,N12892,N12893,N12894,N12895 
	,N12896,N12897,N12898,N12900,N12901,N12902,N12903,N12904 
	,N12905,N12906,N12907,N12908,N12909,N12910,N12912,N12913 
	,N12914,N12915,N12916,N12917,N12918,N12919,N12920,N12921 
	,N12922,N12923,N12924,N12925,N12926,N12927,N12928,N12930 
	,N12931,N12932,N12933,N12934,N12935,N12938,N12939,N12940 
	,N12941,N12942,N12943,N12944,N12945,N12946,N12947,N12948 
	,N12949,N12950,N12951,N12952,N12953,N12955,N12956,N12957 
	,N12958,N12959,N12960,N12961,N12962,N12964,N12965,N12966 
	,N12968,N12969,N12970,N12971,N12972,N12973,N12974,N12975 
	,N12976,N12977,N12978,N12979,N12980,N12981,N12982,N12983 
	,N12984,N12985,N12986,N12987,N12989,N12990,N12991,N12992 
	,N12993,N12994,N12995,N12996,N12997,N12999,N13002,N13003 
	,N13004,N13005,N13006,N13007,N13008,N13009,N13010,N13011 
	,N13012,N13013,N13015,N13016,N13017,N13018,N13019,N13020 
	,N13022,N13023,N13025,N13026,N13027,N13028,N13029,N13031 
	,N13032,N13033,N13034,N13035,N13036,N13037,N13038,N13039 
	,N13040,N13041,N13042,N13043,N13045,N13046,N13047,N13048 
	,N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057 
	,N13058,N13059,N13060,N13061,N13062,N13063,N13064,N13066 
	,N13067,N13068,N13069,N13070,N13071,N13072,N13073,N13074 
	,N13075,N13076,N13077,N13078,N13079,N13080,N13082,N13083 
	,N13084,N13085,N13086,N13088,N13089,N13092,N13093,N13094 
	,N13095,N13096,N13097,N13098,N13099,N13100,N13101,N13102 
	,N13103,N13104,N13105,N13106,N13107,N13108,N13109,N13111 
	,N13112,N13113,N13114,N13115,N13116,N13117,N13119,N13120 
	,N13121,N13122,N13123,N13124,N13125,N13126,N13127,N13128 
	,N13129,N13130,N13131,N13132,N13133,N13134,N13135,N13136 
	,N13137,N13138,N13139,N13140,N13141,N13142,N13143,N13145 
	,N13146,N13147,N13148,N13149,N13150,N13151,N13154,N13155 
	,N13156,N13157,N13158,N13159,N13160,N13161,N13162,N13163 
	,N13164,N13165,N13166,N13167,N13168,N13169,N13170,N13171 
	,N13173,N13174,N13175,N13176,N13177,N13178,N13180,N13181 
	,N13183,N13184,N13185,N13186,N13187,N13188,N13189,N13190 
	,N13191,N13192,N13193,N13195,N13196,N13197,N13198,N13199 
	,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207 
	,N13208,N13209,N13210,N13212,N13213,N13214,N13215,N13216 
	,N13217,N13218,N13219,N13220,N13222,N13223,N13224,N13225 
	,N13227,N13228,N13229,N13230,N13231,N13232,N13233,N13234 
	,N13235,N13236,N13237,N13238,N13239,N13241,N13242,N13243 
	,N13244,N13245,N13247,N13248,N13249,N13251,N13252,N13253 
	,N13254,N13255,N13257,N13258,N13259,N13260,N13261,N13262 
	,N13263,N13264,N13265,N13266,N13267,N13268,N13269,N13270 
	,N13272,N13273,N13274,N13275,N13276,N13277,N13278,N13280 
	,N13281,N13282,N13283,N13284,N13285,N13286,N13287,N13288 
	,N13289,N13290,N13291,N13293,N13295,N13296,N13297,N13298 
	,N13299,N13300,N13301,N13302,N13303,N13304,N13305,N13306 
	,N13307,N13308,N13310,N13311,N13312,N13313,N13314,N13315 
	,N13316,N13317,N13319,N13321,N13322,N13323,N13324,N13325 
	,N13326,N13327,N13328,N13329,N13331,N13332,N13333,N13334 
	,N13335,N13336,N13337,N13339,N13340,N14938,N14940,N14942 
	,N14944,N14945,N14946,N14948,N14949,N14950,N14951,N14954 
	,N14955,N14956,N14957,N14960,N14961,N14963,N14964,N14965 
	,N14966,N14967,N14968,N14970,N14972,N14973,N14974,N14975 
	,N14978,N14979,N14980,N14981,N14982,N14985,N14986,N14988 
	,N14989,N14990,N14991,N14992,N14994,N14995,N14997,N14999 
	,N15000,N15001,N15003,N15006,N15007,N15008,N15009,N15011 
	,N15012,N15013,N15015,N15016,N15017,N15019,N15023,N15024 
	,N15026,N15027,N15028,N15029,N15032,N15033,N15034,N15035 
	,N15036,N15038,N15039,N15041,N15042,N15044,N15047,N15049 
	,N15050,N15051,N15052,N15054,N15055,N15056,N15057,N15061 
	,N15062,N15063,N15064,N15068,N15069,N15071,N15074,N15075 
	,N15076,N15078,N15079,N15081,N15082,N15084,N15086,N15088 
	,N15089,N15090,N15091,N15094,N15096,N15097,N15099,N15100 
	,N15101,N15102,N15103,N15105,N15106,N15107,N15108,N15110 
	,N15111,N15112,N15113,N15114,N15117,N15120,N15121,N15123 
	,N15124,N15125,N15127,N15128,N15129,N15130,N15132,N15133 
	,N15134,N15135,N15136,N15137,N15140,N15141,N15143,N15144 
	,N15145,N15147,N15148,N15150,N15152,N15153,N15154,N15155 
	,N15156,N15159,N15160,N15161,N15162,N15166,N15167,N15168 
	,N15170,N15171,N15172,N15173,N15175,N15176,N15177,N15178 
	,N15181,N15182,N15183,N15184,N15185,N15187,N15188,N15190 
	,N15191,N15192,N15195,N15196,N15199,N15200,N15201,N15202 
	,N15205,N15206,N15207,N15208,N15210,N15211,N15212,N15215 
	,N15216,N15217,N15219,N15221,N15223,N15225,N15226,N15227 
	,N15230,N15231,N15232,N15234,N15235,N15236,N15238,N15239 
	,N15241,N15244,N15246,N15247,N15248,N15249,N15250,N15253 
	,N15254,N15255,N15257,N15260,N15261,N15262,N15263,N15265 
	,N15268,N15270,N15272,N15273,N15274,N15275,N15276,N15278 
	,N15279,N15280,N15281,N15283,N15284,N15286,N15288,N15289 
	,N15290,N15295,N15297,N15298,N15300,N15301,N15302,N15303 
	,N15304,N15306,N15307,N15308,N15309,N15311,N15312,N15313 
	,N15315,N15316,N15317,N15320,N15322,N15323,N15325,N15326 
	,N15327,N15328,N15330,N15331,N15332,N15334,N15335,N15336 
	,N15338,N15339,N15342,N15343,N15345,N15346,N15348,N15349 
	,N15350,N15352,N15353,N15354,N15355,N15356,N15358,N15359 
	,N15360,N15361,N15362,N15363,N15366,N15367,N15369,N15370 
	,N15372,N15373,N15374,N15376,N15377,N15378,N15379,N15380 
	,N15383,N15384,N15385,N15386,N15387,N15390,N15391,N15393 
	,N15394,N15395,N15397,N15399,N15400,N15402,N15403,N15404 
	,N15407,N15408,N15409,N15410,N15412,N15413,N15416,N15417 
	,N15418,N15419,N15420,N15422,N15424,N15426,N15427,N15428 
	,N15429,N15430,N15433,N15434,N15435,N15437,N15440,N15441 
	,N15442,N15444,N15445,N15446,N15448,N15451,N15453,N15455 
	,N15456,N15457,N15458,N15461,N15462,N15463,N15464,N15466 
	,N15467,N15469,N15470,N15471,N15473,N15477,N15479,N15480 
	,N15481,N15482,N15483,N15485,N15487,N15488,N15490,N15492 
	,N15494,N15495,N15496,N15498,N15499,N15503,N15505,N15507 
	,N15508,N15509,N15510,N15511,N15513,N15514,N15515,N15516 
	,N15518,N15519,N15521,N15522,N15523,N15524,N15528,N15530 
	,N15531,N15533,N15534,N15535,N15536,N15539,N15540,N15541 
	,N15543,N15544,N15546,N15547,N15549,N15550,N15553,N15554 
	,N15556,N15557,N15559,N15560,N15561,N15562,N15563,N15565 
	,N15566,N15567,N15568,N15571,N15572,N15573,N15574,N15575 
	,N15578,N15580,N15581,N15583,N15584,N15585,N15587,N15588 
	,N15589,N15590,N15591,N15594,N15595,N15596,N15597,N15598 
	,N15599,N16220,N16294,N16298,N16324,N16328,N16332,N16334 
	,N16343,N16357,N16362,N16376,N16380,N16386,N16390,N16393 
	,N16397,N16401,N16403,N16407,N16409,N16411,N16417,N16464 
	,N16486,N16488,N16489,N16492,N16493,N16494,N16497,N16498 
	,N16500,N16503,N16504,N16505,N16506,N16508,N16509,N16511 
	,N16512,N16514,N16515,N16516,N16517,N16519,N16522,N16523 
	,N16525,N16526,N16528,N16529,N16531,N16533,N16534,N16535 
	,N16537,N16538,N16541,N16542,N16544,N16545,N16546,N16548 
	,N16550,N16551,N16552,N16553,N16554,N16556,N16557,N16558 
	,N16561,N16562,N16564,N16565,N16566,N16567,N16569,N16571 
	,N16636,N16643,N16646,N16662,N16663,N16666,N16667,N16668 
	,N16669,N16673,N16675,N16676,N16677,N16680,N16681,N16682 
	,N16684,N16685,N16686,N16689,N16691,N16692,N16693,N16694 
	,N16697,N16698,N16699,N16703,N16704,N16705,N16708,N16709 
	,N16710,N16711,N16715,N16717,N16718,N16719,N16720,N16722 
	,N16724,N16725,N16726,N16727,N16728,N16731,N16733,N16734 
	,N16737,N16739,N16741,N16742,N16743,N16746,N16748,N16749 
	,N16750,N16752,N16754,N16755,N16756,N16757,N16759,N16761 
	,N16762,N16763,N16764,N16767,N16768,N16769,N16770,N16775 
	,N16776,N16777,N16780,N16781,N16782,N16783,N16786,N16788 
	,N16789,N16790,N16794,N16795,N16796,N16798,N16800,N16801 
	,N16802,N16805,N16808,N16809,N16810,N16811,N16814,N16815 
	,N16816,N16817,N16820,N16822,N16823,N16991,N17141,N17163 
	,N17178,N17198,N17202,N17205,N17207,N17211,N17213,N17217 
	,N17220,N17223,N17227,N17230,N17234,N17237,N17239,N17244 
	,N17247,N17251,N17254,N17256,N17263,N17267,N17270,N23218 
	,N23226,N23239,N23240,N23255,N23273,N23274,N23275,N23276 
	,N23277,N23278,N23282,N23285,N23286,N23288,N23290,N23296 
	,N23302,N23303,N23304,N23307,N23308,N23309,N23312,N23313 
	,N23314,N23315,N23318,N23319,N23320,N23321,N23322,N23324 
	,N23344,N23358,N23367,N23375,N23383,N23391,N23399,N23407 
	,N23415,N23421,N23433,N23439,N23456,N44729,N44730,N44974 
	,N44981,N44986,N45000,N45002,N45015,N45016,N45019,N45020 
	,N45023,N45025,N45027,N45031,N45032,N45033,N45036,N45040 
	,N45043,N45045,N45046,N45050,N45051,N45052,N45055,N45061 
	,N45064,N45065,N45067,N45068,N45070,N45071,N45072,N45115 
	,N45117,N45118,N45119,N45122,N45128,N45132,N45139,N45146 
	,N45148,N45150,N45152,N45155,N45159,N45190,N45195,N45200 
	,N45203,N45206,N45208,N45238,N45239,N45242,N45245,N45246 
	,N45249,N45252,N45254,N45259,N45262,N45267,N45270,N45273 
	,N45276,N45279,N45282,N45283,N45286,N45290,N45293,N45296 
	,N45297,N45300,N45341,N45342,N45345,N45350,N45353,N45355 
	,N45358,N45368,N45371,N45377,N45380,N45383,N45386,N45389 
	,N45391,N45394,N45397,N45400,N45439,N45446,N45451,N45454 
	,N45456,N45460,N45464,N45473,N45494,N45499,N45504,N45518 
	,N45525,N45526,N45530,N45533,N45547,N45549,N45552,N45569 
	,N45572,N45575,N45576,N45581,N45583,N45584,N45587,N45592 
	,N45595,N45598,N45601,N45604,N45608,N45611,N45612,N45615 
	,N45618,N45620,N45621,N45624,N45631,N45668,N45677,N45679 
	,N45684,N45687,N45692,N45695,N45698,N45700,N45705,N45708 
	,N45711,N45713,N45718,N45720,N45721,N45724,N45756,N45763 
	,N45771,N45774,N45780,N45786,N45792,N45799,N45805,N45811 
	,N45817,N45823,N45829,N45835,N45841,N45847,N45854;
INVX2 inst_blk01_cellmath__39_I509 (.Y(N5740), .A(a_man[0]));
CLKINVX12 inst_blk01_cellmath__39_I510 (.Y(N5723), .A(a_man[1]));
CLKINVX6 inst_blk01_cellmath__39_I511 (.Y(N6122), .A(a_man[2]));
INVX3 inst_blk01_cellmath__39_I512 (.Y(N5716), .A(a_man[3]));
CLKINVX6 inst_blk01_cellmath__39_I513 (.Y(N5995), .A(a_man[4]));
CLKINVX6 inst_blk01_cellmath__39_I514 (.Y(N6378), .A(a_man[5]));
INVX12 inst_blk01_cellmath__39_I515 (.Y(N5927), .A(a_man[6]));
CLKINVX6 inst_blk01_cellmath__39_I516 (.Y(N6263), .A(a_man[7]));
CLKINVX4 inst_blk01_cellmath__39_I517 (.Y(N5778), .A(a_man[8]));
CLKINVX6 inst_blk01_cellmath__39_I518 (.Y(N6155), .A(a_man[9]));
CLKINVX8 inst_blk01_cellmath__39_I519 (.Y(N5662), .A(a_man[10]));
INVX2 inst_blk01_cellmath__39_I520 (.Y(N6041), .A(a_man[11]));
INVX3 inst_blk01_cellmath__39_I521 (.Y(N5565), .A(a_man[12]));
CLKINVX8 inst_blk01_cellmath__39_I522 (.Y(N5929), .A(a_man[13]));
CLKINVX4 inst_blk01_cellmath__39_I523 (.Y(N6308), .A(a_man[14]));
INVX2 inst_blk01_cellmath__39_I524 (.Y(N5821), .A(a_man[15]));
INVX3 inst_blk01_cellmath__39_I526 (.Y(N6201), .A(a_man[16]));
INVX3 inst_blk01_cellmath__39_I527 (.Y(N5705), .A(a_man[17]));
INVX2 inst_blk01_cellmath__39_I528 (.Y(N6089), .A(a_man[18]));
INVX2 inst_blk01_cellmath__39_I529 (.Y(N5605), .A(a_man[19]));
INVX1 inst_blk01_cellmath__39_I530 (.Y(N5981), .A(a_man[20]));
BUFX3 inst_blk01_cellmath__39_I531 (.Y(N5637), .A(N5981));
INVX2 inst_blk01_cellmath__39_I532 (.Y(N6354), .A(a_man[21]));
INVX1 inst_blk01_cellmath__39_I533 (.Y(N5870), .A(a_man[22]));
BUFX2 inst_blk01_cellmath__39_I534 (.Y(N6010), .A(N5870));
XNOR2X1 inst_blk01_cellmath__39_I535 (.Y(N5980), .A(a_man[9]), .B(a_man[2]));
OR2XL inst_blk01_cellmath__39_I536 (.Y(N6171), .A(a_man[9]), .B(a_man[2]));
ADDFX1 inst_blk01_cellmath__39_I537 (.CO(N6056), .S(N5872), .A(a_man[3]), .B(a_man[10]), .CI(N5723));
ADDFXL inst_blk01_cellmath__39_I538 (.CO(N5578), .S(N6246), .A(N6122), .B(a_man[11]), .CI(a_man[4]));
ADDFXL inst_blk01_cellmath__39_I539 (.CO(N5947), .S(N5755), .A(a_man[5]), .B(a_man[12]), .CI(N5716));
ADDFX1 inst_blk01_cellmath__39_I540 (.CO(N6322), .S(N6136), .A(a_man[6]), .B(a_man[13]), .CI(N5995));
XNOR2X1 inst_blk01_cellmath__39_I541 (.Y(N5650), .A(a_man[14]), .B(a_man[7]));
OR2XL inst_blk01_cellmath__39_I542 (.Y(N5839), .A(a_man[14]), .B(a_man[7]));
OR2XL inst_blk01_cellmath__39_I545 (.Y(N6105), .A(a_man[15]), .B(a_man[8]));
OR2XL inst_blk01_cellmath__39_I548 (.Y(N6374), .A(a_man[16]), .B(a_man[9]));
XNOR2X1 inst_blk01_cellmath__39_I551 (.Y(N5960), .A(a_man[17]), .B(a_man[10]));
OR2XL inst_blk01_cellmath__39_I552 (.Y(N6152), .A(a_man[17]), .B(a_man[10]));
ADDFXL inst_blk01_cellmath__39_I553 (.CO(N6038), .S(N5854), .A(N5778), .B(a_man[1]), .CI(N5716));
ADDHX1 inst_blk01_cellmath__39_I554 (.CO(N5562), .S(N6225), .A(N5565), .B(N5981));
ADDFX1 inst_blk01_cellmath__39_I555 (.CO(N5925), .S(N5736), .A(a_man[11]), .B(a_man[18]), .CI(a_man[2]));
ADDFHXL inst_blk01_cellmath__39_I556 (.CO(N6305), .S(N6120), .A(N5995), .B(N5929), .CI(N6155));
XNOR2X1 inst_blk01_cellmath__39_I557 (.Y(N5629), .A(a_man[19]), .B(a_man[12]));
OR2XL inst_blk01_cellmath__39_I558 (.Y(N5819), .A(a_man[19]), .B(a_man[12]));
ADDFHXL inst_blk01_cellmath__39_I559 (.CO(N5702), .S(N6391), .A(a_man[3]), .B(a_man[0]), .CI(N6378));
ADDHX1 inst_blk01_cellmath__39_I560 (.CO(N6087), .S(N5896), .A(N5662), .B(N6308));
XNOR2X1 inst_blk01_cellmath__39_I561 (.Y(N6276), .A(a_man[20]), .B(a_man[13]));
OR2XL inst_blk01_cellmath__39_I562 (.Y(N5601), .A(a_man[20]), .B(a_man[13]));
ADDFX1 inst_blk01_cellmath__39_I563 (.CO(N6351), .S(N6167), .A(a_man[4]), .B(a_man[1]), .CI(N5927));
ADDHX1 inst_blk01_cellmath__39_I564 (.CO(N5867), .S(N5674), .A(N6041), .B(N5821));
ADDFHX1 inst_blk01_cellmath__39_I565 (.CO(N6243), .S(N6054), .A(a_man[14]), .B(a_man[21]), .CI(a_man[0]));
ADDFHXL inst_blk01_cellmath__39_I566 (.CO(N5752), .S(N5574), .A(a_man[5]), .B(a_man[2]), .CI(N6263));
ADDHX1 inst_blk01_cellmath__39_I567 (.CO(N6133), .S(N5942), .A(N5565), .B(N6201));
XNOR2X1 inst_blk01_cellmath__39_I568 (.Y(N6318), .A(a_man[22]), .B(a_man[15]));
OR2XL inst_blk01_cellmath__39_I569 (.Y(N5646), .A(a_man[22]), .B(a_man[15]));
ADDFX1 inst_blk01_cellmath__39_I570 (.CO(N6407), .S(N6214), .A(a_man[3]), .B(a_man[1]), .CI(a_man[6]));
ADDFXL inst_blk01_cellmath__39_I571 (.CO(N5910), .S(N5717), .A(N5778), .B(N5705), .CI(N5929));
ADDFXL inst_blk01_cellmath__39_I572 (.CO(N6289), .S(N6101), .A(a_man[2]), .B(a_man[16]), .CI(a_man[4]));
ADDFXL inst_blk01_cellmath__39_I573 (.CO(N5803), .S(N5616), .A(a_man[7]), .B(N6308), .CI(N6155));
ADDFX1 inst_blk01_cellmath__39_I574 (.CO(N6182), .S(N5988), .A(a_man[3]), .B(a_man[17]), .CI(a_man[5]));
ADDHX1 inst_blk01_cellmath__39_I575 (.CO(N5686), .S(N6370), .A(N5662), .B(a_man[8]));
ADDFX1 inst_blk01_cellmath__39_I576 (.CO(N6070), .S(N5883), .A(a_man[4]), .B(a_man[18]), .CI(a_man[6]));
ADDHX1 inst_blk01_cellmath__39_I577 (.CO(N5589), .S(N6255), .A(a_man[9]), .B(N6041));
ADDFX1 inst_blk01_cellmath__39_I578 (.CO(N5956), .S(N5769), .A(a_man[5]), .B(a_man[19]), .CI(a_man[7]));
ADDHX1 inst_blk01_cellmath__39_I579 (.CO(N6336), .S(N6148), .A(a_man[10]), .B(N5565));
ADDFX1 inst_blk01_cellmath__39_I580 (.CO(N5849), .S(N5656), .A(a_man[6]), .B(a_man[20]), .CI(a_man[8]));
ADDHX1 inst_blk01_cellmath__39_I581 (.CO(N6223), .S(N6034), .A(N5929), .B(a_man[11]));
ADDFXL inst_blk01_cellmath__39_I582 (.CO(N5732), .S(N6421), .A(a_man[7]), .B(a_man[21]), .CI(a_man[9]));
XNOR2X1 inst_blk01_cellmath__39_I583 (.Y(N5922), .A(a_man[22]), .B(a_man[8]));
OR2XL inst_blk01_cellmath__39_I584 (.Y(N6115), .A(a_man[22]), .B(a_man[8]));
XNOR2X1 inst_blk01_cellmath__39_I585 (.Y(N5815), .A(a_man[5]), .B(N5740));
OR2XL inst_blk01_cellmath__39_I586 (.Y(N6002), .A(a_man[5]), .B(N5740));
ADDFX1 inst_blk01_cellmath__39_I587 (.CO(N5894), .S(N5699), .A(N5723), .B(a_man[6]), .CI(N5821));
ADDFX1 inst_blk01_cellmath__39_I588 (.CO(N6272), .S(N6084), .A(a_man[0]), .B(a_man[7]), .CI(N6122));
ADDHX1 inst_blk01_cellmath__39_I589 (.CO(N5786), .S(N5598), .A(N5929), .B(N6201));
ADDFX1 inst_blk01_cellmath__39_I590 (.CO(N6163), .S(N5971), .A(a_man[1]), .B(a_man[8]), .CI(N5716));
ADDFX1 inst_blk01_cellmath__39_I591 (.CO(N5669), .S(N6347), .A(N5705), .B(N6041), .CI(N6308));
ADDFX1 inst_blk01_cellmath__39_I592 (.CO(N6050), .S(N5862), .A(N5740), .B(N6089), .CI(N5995));
ADDFX1 inst_blk01_cellmath__39_I593 (.CO(N5570), .S(N6237), .A(N5565), .B(N5821), .CI(N5980));
ADDFX1 inst_blk01_cellmath__39_I594 (.CO(N5937), .S(N5748), .A(N6201), .B(N6378), .CI(N5605));
ADDFX1 inst_blk01_cellmath__39_I595 (.CO(N6314), .S(N6127), .A(N6171), .B(N5929), .CI(N5872));
ADDFXL inst_blk01_cellmath__39_I596 (.CO(N5828), .S(N5640), .A(N5637), .B(N5705), .CI(N5927));
ADDFX1 inst_blk01_cellmath__39_I597 (.CO(N6207), .S(N6013), .A(N6056), .B(N6308), .CI(N6246));
ADDFX1 inst_blk01_cellmath__39_I598 (.CO(N5713), .S(N6399), .A(N6354), .B(N6089), .CI(N6263));
ADDFX1 inst_blk01_cellmath__39_I599 (.CO(N6096), .S(N5906), .A(N5578), .B(N5821), .CI(N5755));
ADDHX1 inst_blk01_cellmath__39_I29553 (.CO(N5776), .S(N45273), .A(N5870), .B(N6041));
ADDFX1 inst_blk01_cellmath__39_I29552 (.CO(N6259), .S(N45245), .A(a_man[0]), .B(N6122), .CI(N6263));
ADDFXL inst_blk01_cellmath__39_I608 (.CO(N6030), .S(N5843), .A(N5776), .B(N6374), .CI(N6259));
ADDFXL inst_blk01_cellmath__39_I609 (.CO(N6416), .S(N6220), .A(N5960), .B(N6225), .CI(N5854));
ADDFX1 inst_blk01_cellmath__39_I610 (.CO(N5918), .S(N5727), .A(N6152), .B(N6354), .CI(N5562));
ADDFX1 inst_blk01_cellmath__39_I611 (.CO(N6297), .S(N6110), .A(N6038), .B(N6120), .CI(N5736));
ADDFHXL inst_blk01_cellmath__39_I612 (.CO(N5810), .S(N5623), .A(N5925), .B(N6010), .CI(N6305));
ADDFHXL inst_blk01_cellmath__39_I613 (.CO(N6192), .S(N5998), .A(N5896), .B(N5629), .CI(N6391));
ADDFX1 inst_blk01_cellmath__39_I614 (.CO(N5695), .S(N6381), .A(N6087), .B(N5819), .CI(N5702));
ADDFX1 inst_blk01_cellmath__39_I615 (.CO(N6079), .S(N5891), .A(N6276), .B(N5674), .CI(N6167));
ADDFXL inst_blk01_cellmath__39_I616 (.CO(N5595), .S(N6267), .A(N5601), .B(N5867), .CI(N6351));
ADDFX1 inst_blk01_cellmath__39_I617 (.CO(N5966), .S(N5780), .A(N6054), .B(N5942), .CI(N5574));
ADDFHXL inst_blk01_cellmath__39_I618 (.CO(N6343), .S(N6157), .A(N6133), .B(N6243), .CI(N5752));
ADDFX1 inst_blk01_cellmath__39_I619 (.CO(N5857), .S(N5664), .A(N6318), .B(N6214), .CI(N5717));
ADDFX1 inst_blk01_cellmath__39_I620 (.CO(N6233), .S(N6045), .A(N5646), .B(N6089), .CI(N6407));
ADDFXL inst_blk01_cellmath__39_I621 (.CO(N5742), .S(N5566), .A(N5910), .B(N6101), .CI(N5616));
ADDFXL inst_blk01_cellmath__39_I622 (.CO(N6123), .S(N5933), .A(N5605), .B(N5821), .CI(N6289));
ADDFX1 inst_blk01_cellmath__39_I623 (.CO(N5635), .S(N6310), .A(N5803), .B(N6370), .CI(N5988));
ADDFX1 inst_blk01_cellmath__39_I624 (.CO(N6009), .S(N5824), .A(N5637), .B(N5686), .CI(N6201));
ADDFX1 inst_blk01_cellmath__39_I625 (.CO(N6396), .S(N6204), .A(N6182), .B(N6255), .CI(N5883));
ADDFX1 inst_blk01_cellmath__39_I626 (.CO(N5903), .S(N5708), .A(N6354), .B(N5705), .CI(N5589));
ADDFX1 inst_blk01_cellmath__39_I627 (.CO(N6281), .S(N6092), .A(N6070), .B(N6148), .CI(N5769));
ADDFX1 inst_blk01_cellmath__39_I628 (.CO(N5793), .S(N5609), .A(N6010), .B(N6089), .CI(N6336));
ADDFXL inst_blk01_cellmath__39_I629 (.CO(N6174), .S(N5983), .A(N6034), .B(N5956), .CI(N5656));
ADDFX1 inst_blk01_cellmath__39_I630 (.CO(N5680), .S(N6357), .A(N5605), .B(a_man[12]), .CI(N6308));
ADDFX1 inst_blk01_cellmath__39_I631 (.CO(N6060), .S(N5876), .A(N5849), .B(N6223), .CI(N6421));
ADDFX1 inst_blk01_cellmath__39_I632 (.CO(N5581), .S(N6248), .A(a_man[13]), .B(a_man[10]), .CI(N5821));
ADDFX1 inst_blk01_cellmath__39_I633 (.CO(N5949), .S(N5759), .A(N5637), .B(N5732), .CI(N5922));
ADDFX1 inst_blk01_cellmath__39_I634 (.CO(N6326), .S(N6141), .A(a_man[11]), .B(a_man[9]), .CI(a_man[14]));
ADDFX1 inst_blk01_cellmath__39_I635 (.CO(N5840), .S(N5651), .A(N6115), .B(N6354), .CI(N6201));
ADDFX1 inst_blk01_cellmath__39_I636 (.CO(N6218), .S(N6025), .A(a_man[12]), .B(a_man[10]), .CI(a_man[15]));
ADDHX1 inst_blk01_cellmath__39_I637 (.CO(N5721), .S(N6413), .A(N5705), .B(N6010));
ADDFX1 inst_blk01_cellmath__39_I638 (.CO(N6108), .S(N5915), .A(a_man[13]), .B(a_man[11]), .CI(a_man[16]));
XNOR2X1 inst_blk01_cellmath__39_I639 (.Y(N6292), .A(a_man[12]), .B(a_man[14]));
OR2XL inst_blk01_cellmath__39_I640 (.Y(N5621), .A(a_man[12]), .B(a_man[14]));
XNOR2X1 inst_blk01_cellmath__39_I641 (.Y(N6190), .A(a_man[13]), .B(a_man[15]));
OR2XL inst_blk01_cellmath__39_I642 (.Y(N6377), .A(a_man[13]), .B(a_man[15]));
XNOR2X1 inst_blk01_cellmath__39_I643 (.Y(N6077), .A(a_man[14]), .B(a_man[16]));
OR2XL inst_blk01_cellmath__39_I644 (.Y(N6261), .A(a_man[14]), .B(a_man[16]));
XNOR2X1 inst_blk01_cellmath__39_I645 (.Y(N5962), .A(a_man[15]), .B(a_man[17]));
OR2XL inst_blk01_cellmath__39_I646 (.Y(N6154), .A(a_man[15]), .B(a_man[17]));
INVXL inst_blk01_cellmath__39_I647 (.Y(N5739), .A(N5927));
ADDHX1 inst_blk01_cellmath__39_I648 (.CO(N5820), .S(N5631), .A(N5995), .B(N6263));
ADDHX1 inst_blk01_cellmath__39_I649 (.CO(N6200), .S(N6007), .A(N6378), .B(N5778));
ADDFX1 inst_blk01_cellmath__39_I650 (.CO(N5703), .S(N6392), .A(N6155), .B(a_man[0]), .CI(N5927));
ADDFX1 inst_blk01_cellmath__39_I651 (.CO(N6088), .S(N5899), .A(N5662), .B(a_man[1]), .CI(N6263));
ADDFX1 inst_blk01_cellmath__39_I652 (.CO(N5604), .S(N6278), .A(N6041), .B(a_man[2]), .CI(N5778));
ADDFX1 inst_blk01_cellmath__39_I653 (.CO(N5976), .S(N5789), .A(a_man[3]), .B(N5565), .CI(N6155));
ADDFX1 inst_blk01_cellmath__39_I654 (.CO(N6352), .S(N6169), .A(N5929), .B(a_man[4]), .CI(N5662));
ADDFX1 inst_blk01_cellmath__39_I655 (.CO(N5869), .S(N5675), .A(N6308), .B(N5778), .CI(N6041));
ADDFX1 inst_blk01_cellmath__39_I656 (.CO(N6244), .S(N6055), .A(N6002), .B(N5565), .CI(N6155));
ADDFX1 inst_blk01_cellmath__39_I657 (.CO(N5754), .S(N5575), .A(N5894), .B(N5598), .CI(N5662));
ADDFXL inst_blk01_cellmath__39_I658 (.CO(N6134), .S(N5945), .A(N6272), .B(N5786), .CI(N5971));
ADDFX1 inst_blk01_cellmath__39_I659 (.CO(N5648), .S(N6320), .A(N5669), .B(N6163), .CI(N5862));
ADDFX1 inst_blk01_cellmath__39_I660 (.CO(N6021), .S(N5837), .A(N5748), .B(N6050), .CI(N5570));
ADDFXL inst_blk01_cellmath__39_I661 (.CO(N6409), .S(N6215), .A(N5640), .B(N5937), .CI(N6314));
ADDFHXL inst_blk01_cellmath__39_I662 (.CO(N5911), .S(N5718), .A(N5828), .B(N6399), .CI(N6207));
ADDFX1 inst_blk01_cellmath__39_I29554 (.CO(N45252), .S(N6285), .A(N5778), .B(N5605), .CI(N6010));
ADDFXL inst_blk01_cellmath__39_I663 (.CO(N6290), .S(N6103), .A(N6285), .B(N5713), .CI(N6096));
ADDFHXL inst_blk01_cellmath__39_I29550 (.CO(N45282), .S(N45267), .A(N5927), .B(N5723), .CI(N5662));
ADDFHXL inst_blk01_cellmath__39_I29560 (.CO(N6144), .S(N45276), .A(N6105), .B(N5605), .CI(N45282));
XNOR2X1 inst_blk01_cellmath__39_I29551 (.Y(N45296), .A(a_man[16]), .B(a_man[9]));
ADDFX1 inst_blk01_cellmath__39_I29561 (.CO(N5653), .S(N45239), .A(N45296), .B(N45273), .CI(N45245));
ADDFHXL inst_blk01_cellmath__39_I667 (.CO(N6072), .S(N5885), .A(N5843), .B(N6144), .CI(N5653));
ADDFXL inst_blk01_cellmath__39_I668 (.CO(N5591), .S(N6256), .A(N5727), .B(N6030), .CI(N6416));
ADDFXL inst_blk01_cellmath__39_I669 (.CO(N5958), .S(N5774), .A(N5623), .B(N5918), .CI(N6297));
ADDFHXL inst_blk01_cellmath__39_I670 (.CO(N6337), .S(N6150), .A(N5810), .B(N6192), .CI(N6381));
ADDFXL inst_blk01_cellmath__39_I671 (.CO(N5852), .S(N5659), .A(N6267), .B(N5695), .CI(N6079));
ADDFXL inst_blk01_cellmath__39_I672 (.CO(N6224), .S(N6036), .A(N5595), .B(N6157), .CI(N5966));
ADDFHXL inst_blk01_cellmath__39_I673 (.CO(N5734), .S(N5560), .A(N6343), .B(N6045), .CI(N5857));
ADDFXL inst_blk01_cellmath__39_I674 (.CO(N6117), .S(N5923), .A(N5933), .B(N6233), .CI(N5742));
ADDFXL inst_blk01_cellmath__39_I675 (.CO(N5627), .S(N6303), .A(N5824), .B(N6123), .CI(N5635));
ADDFHXL inst_blk01_cellmath__39_I676 (.CO(N6004), .S(N5817), .A(N5708), .B(N6009), .CI(N6396));
ADDFHXL inst_blk01_cellmath__39_I677 (.CO(N6388), .S(N6197), .A(N5609), .B(N5903), .CI(N6281));
ADDFXL inst_blk01_cellmath__39_I678 (.CO(N5895), .S(N5700), .A(N5793), .B(N6357), .CI(N6174));
ADDFXL inst_blk01_cellmath__39_I679 (.CO(N6274), .S(N6085), .A(N6248), .B(N5680), .CI(N6060));
ADDFX1 inst_blk01_cellmath__39_I680 (.CO(N5787), .S(N5600), .A(N6141), .B(N5581), .CI(N5949));
ADDFX1 inst_blk01_cellmath__39_I681 (.CO(N6166), .S(N5973), .A(N6025), .B(N6326), .CI(N6413));
ADDFX1 inst_blk01_cellmath__39_I682 (.CO(N5671), .S(N6348), .A(N6089), .B(N6218), .CI(N5721));
ADDFX1 inst_blk01_cellmath__39_I683 (.CO(N6051), .S(N5866), .A(a_man[17]), .B(N6108), .CI(N5605));
ADDFX1 inst_blk01_cellmath__39_I684 (.CO(N5572), .S(N6241), .A(N5637), .B(a_man[18]), .CI(N5621));
ADDFX1 inst_blk01_cellmath__39_I685 (.CO(N5940), .S(N5749), .A(N6354), .B(a_man[19]), .CI(N6377));
ADDFX1 inst_blk01_cellmath__39_I686 (.CO(N6317), .S(N6131), .A(N6010), .B(a_man[20]), .CI(N6261));
ADDFX1 inst_blk01_cellmath__39_I687 (.CO(N5833), .S(N5644), .A(a_man[21]), .B(a_man[18]), .CI(N6201));
ADDFX1 inst_blk01_cellmath__39_I688 (.CO(N6212), .S(N6017), .A(a_man[19]), .B(a_man[17]), .CI(a_man[22]));
INVXL inst_blk01_cellmath__39_I689 (.Y(N6405), .A(N5716));
ADDHXL inst_blk01_cellmath__39_I690 (.CO(N5615), .S(N6288), .A(N5723), .B(N5995));
ADDHX1 inst_blk01_cellmath__39_I691 (.CO(N5987), .S(N5802), .A(N6378), .B(N6122));
ADDFX1 inst_blk01_cellmath__39_I692 (.CO(N6369), .S(N6180), .A(N5739), .B(N5740), .CI(N5716));
ADDFXL inst_blk01_cellmath__39_I693 (.CO(N5882), .S(N5685), .A(N5723), .B(N5631), .CI(N5927));
ADDFX1 inst_blk01_cellmath__39_I694 (.CO(N6254), .S(N6069), .A(N5820), .B(N6122), .CI(N6007));
ADDFX1 inst_blk01_cellmath__39_I695 (.CO(N5767), .S(N5588), .A(N6200), .B(N6392), .CI(N5716));
ADDFX1 inst_blk01_cellmath__39_I696 (.CO(N6147), .S(N5954), .A(N5703), .B(N5899), .CI(N5995));
ADDFX1 inst_blk01_cellmath__39_I697 (.CO(N5655), .S(N6335), .A(N6278), .B(N6088), .CI(N6378));
ADDFXL inst_blk01_cellmath__39_I698 (.CO(N6033), .S(N5847), .A(N5789), .B(N5604), .CI(N5927));
ADDFX1 inst_blk01_cellmath__39_I699 (.CO(N6419), .S(N6222), .A(N6169), .B(N5976), .CI(N6263));
ADDFX1 inst_blk01_cellmath__39_I700 (.CO(N5921), .S(N5730), .A(N5815), .B(N6352), .CI(N5675));
ADDFX1 inst_blk01_cellmath__39_I701 (.CO(N6301), .S(N6114), .A(N5699), .B(N5869), .CI(N6055));
ADDFX1 inst_blk01_cellmath__39_I702 (.CO(N5813), .S(N5626), .A(N6244), .B(N6084), .CI(N5575));
ADDFX1 inst_blk01_cellmath__39_I703 (.CO(N6194), .S(N6001), .A(N5754), .B(N6347), .CI(N5945));
ADDFX1 inst_blk01_cellmath__39_I704 (.CO(N5698), .S(N6385), .A(N6237), .B(N6134), .CI(N6320));
ADDFXL inst_blk01_cellmath__39_I705 (.CO(N6082), .S(N5893), .A(N6127), .B(N5837), .CI(N5648));
ADDFXL inst_blk01_cellmath__39_I706 (.CO(N5597), .S(N6270), .A(N6021), .B(N6013), .CI(N6215));
ADDFHXL inst_blk01_cellmath__39_I707 (.CO(N5969), .S(N5785), .A(N5906), .B(N6409), .CI(N5718));
ADDFHXL inst_blk01_cellmath__39_I29555 (.CO(N45279), .S(N5799), .A(N5947), .B(N6201), .CI(N6136));
ADDFX1 inst_blk01_cellmath__39_I708 (.CO(N6346), .S(N6162), .A(N5911), .B(N5799), .CI(N6103));
ADDHX1 inst_blk01_cellmath__39_I29548 (.CO(N45238), .S(N45290), .A(N6378), .B(N5740));
ADDFX1 inst_blk01_cellmath__39_I29557 (.CO(N45270), .S(N5683), .A(N6322), .B(N5650), .CI(N45290));
ADDFX1 inst_blk01_cellmath__39_I29556 (.CO(N45242), .S(N45293), .A(N5705), .B(N5637), .CI(N6155));
ADDFHXL inst_blk01_cellmath__39_I29562 (.CO(N45283), .S(N5618), .A(N45293), .B(N45252), .CI(N45279));
ADDFHX1 inst_blk01_cellmath__39_I709 (.CO(N5861), .S(N5668), .A(N5683), .B(N6290), .CI(N5618));
ADDFX1 inst_blk01_cellmath__39_I29558 (.CO(N45300), .S(N45286), .A(N6089), .B(N6354), .CI(N5839));
XNOR2X1 inst_blk01_cellmath__39_I29549 (.Y(N45254), .A(a_man[15]), .B(a_man[8]));
ADDFHXL inst_blk01_cellmath__39_I29559 (.CO(N45262), .S(N45249), .A(N45254), .B(N45238), .CI(N45267));
ADDFHXL inst_blk01_cellmath__39_I29564 (.CO(N5687), .S(N45259), .A(N45300), .B(N45276), .CI(N45262));
ADDFHXL inst_blk01_cellmath__39_I712 (.CO(N6126), .S(N5935), .A(N5687), .B(N6220), .CI(N5885));
ADDFHX1 inst_blk01_cellmath__39_I713 (.CO(N5638), .S(N6313), .A(N6072), .B(N6110), .CI(N6256));
ADDFXL inst_blk01_cellmath__39_I714 (.CO(N6012), .S(N5827), .A(N5998), .B(N5591), .CI(N5774));
ADDFHXL inst_blk01_cellmath__39_I715 (.CO(N6398), .S(N6206), .A(N5958), .B(N5891), .CI(N6150));
ADDFXL inst_blk01_cellmath__39_I716 (.CO(N5905), .S(N5710), .A(N6337), .B(N5780), .CI(N5659));
ADDFHX1 inst_blk01_cellmath__39_I717 (.CO(N6284), .S(N6095), .A(N5852), .B(N5664), .CI(N6036));
ADDFHX1 inst_blk01_cellmath__39_I718 (.CO(N5798), .S(N5611), .A(N6224), .B(N5566), .CI(N5560));
ADDFHX1 inst_blk01_cellmath__39_I719 (.CO(N6175), .S(N5984), .A(N6310), .B(N5734), .CI(N5923));
ADDFHX1 inst_blk01_cellmath__39_I720 (.CO(N5682), .S(N6363), .A(N6117), .B(N6204), .CI(N6303));
ADDFHX1 inst_blk01_cellmath__39_I721 (.CO(N6064), .S(N5878), .A(N5627), .B(N6092), .CI(N5817));
ADDFHX1 inst_blk01_cellmath__39_I722 (.CO(N5582), .S(N6250), .A(N6004), .B(N5983), .CI(N6197));
ADDFHXL inst_blk01_cellmath__39_I723 (.CO(N5950), .S(N5763), .A(N6388), .B(N5876), .CI(N5700));
ADDFHXL inst_blk01_cellmath__39_I724 (.CO(N6330), .S(N6142), .A(N5895), .B(N5759), .CI(N6085));
ADDFXL inst_blk01_cellmath__39_I725 (.CO(N5842), .S(N5652), .A(N6274), .B(N5651), .CI(N5600));
ADDFX1 inst_blk01_cellmath__39_I726 (.CO(N6219), .S(N6029), .A(N5973), .B(N5840), .CI(N5787));
ADDFX1 inst_blk01_cellmath__39_I727 (.CO(N5725), .S(N6414), .A(N6348), .B(N5915), .CI(N6166));
ADDFX1 inst_blk01_cellmath__39_I728 (.CO(N6109), .S(N5916), .A(N5671), .B(N6292), .CI(N5866));
ADDFX1 inst_blk01_cellmath__39_I729 (.CO(N5622), .S(N6296), .A(N6051), .B(N6190), .CI(N6241));
ADDFX1 inst_blk01_cellmath__39_I730 (.CO(N5997), .S(N5808), .A(N5572), .B(N6077), .CI(N5749));
ADDFX1 inst_blk01_cellmath__39_I731 (.CO(N6379), .S(N6191), .A(N5940), .B(N5962), .CI(N6131));
ADDFX1 inst_blk01_cellmath__39_I732 (.CO(N5889), .S(N5693), .A(N5644), .B(N6154), .CI(N6317));
ADDFX1 inst_blk01_cellmath__39_I733 (.CO(N6266), .S(N6078), .A(N5833), .B(a_man[16]), .CI(N6017));
ADDFX1 inst_blk01_cellmath__39_I734 (.CO(N5779), .S(N5594), .A(a_man[20]), .B(a_man[18]), .CI(N6212));
ADDHX1 inst_blk01_cellmath__39_I735 (.CO(N6156), .S(N5965), .A(a_man[19]), .B(a_man[21]));
ADDHX1 inst_blk01_cellmath__39_I736 (.CO(N5663), .S(N6341), .A(a_man[20]), .B(a_man[22]));
NOR2XL inst_blk01_cellmath__39_I739 (.Y(N6309), .A(N6405), .B(N5740));
NAND2XL inst_blk01_cellmath__39_I740 (.Y(N5634), .A(N5740), .B(N6405));
NOR2XL inst_blk01_cellmath__39_I741 (.Y(N5823), .A(N5716), .B(N6288));
NOR2XL inst_blk01_cellmath__39_I743 (.Y(N6203), .A(N5615), .B(N5802));
NAND2XL inst_blk01_cellmath__39_I744 (.Y(N6395), .A(N5615), .B(N5802));
NOR2XL inst_blk01_cellmath__39_I745 (.Y(N5706), .A(N5987), .B(N6180));
NAND2XL inst_blk01_cellmath__39_I746 (.Y(N5901), .A(N5987), .B(N6180));
NOR2X1 inst_blk01_cellmath__39_I747 (.Y(N6091), .A(N6369), .B(N5685));
NOR2XL inst_blk01_cellmath__39_I749 (.Y(N5607), .A(N5882), .B(N6069));
NAND2X1 inst_blk01_cellmath__39_I750 (.Y(N5792), .A(N5882), .B(N6069));
NOR2XL inst_blk01_cellmath__39_I751 (.Y(N5982), .A(N6254), .B(N5588));
NAND2XL inst_blk01_cellmath__39_I752 (.Y(N6173), .A(N6254), .B(N5588));
NOR2XL inst_blk01_cellmath__39_I753 (.Y(N6356), .A(N5767), .B(N5954));
NAND2XL inst_blk01_cellmath__39_I754 (.Y(N5677), .A(N5767), .B(N5954));
NOR2XL inst_blk01_cellmath__39_I755 (.Y(N5875), .A(N6147), .B(N6335));
NOR2XL inst_blk01_cellmath__39_I757 (.Y(N6247), .A(N5655), .B(N5847));
NAND2XL inst_blk01_cellmath__39_I758 (.Y(N5580), .A(N5655), .B(N5847));
NOR2XL inst_blk01_cellmath__39_I759 (.Y(N5758), .A(N6033), .B(N6222));
NOR2XL inst_blk01_cellmath__39_I761 (.Y(N6138), .A(N6419), .B(N5730));
NAND2XL inst_blk01_cellmath__39_I762 (.Y(N6325), .A(N6419), .B(N5730));
NAND3XL inst_blk01_cellmath__39_I10659 (.Y(N6188), .A(N5723), .B(N6122), .C(N5740));
AOI21XL inst_blk01_cellmath__39_I765 (.Y(N6339), .A0(N5634), .A1(N6188), .B0(N6309));
AOI21XL inst_blk01_cellmath__39_I766 (.Y(N6227), .A0(N6395), .A1(N5823), .B0(N6203));
OAI2BB1X1 inst_blk01_cellmath__39_I10660 (.Y(N5563), .A0N(N5716), .A1N(N6288), .B0(N6395));
OAI21XL inst_blk01_cellmath__39_I768 (.Y(N5898), .A0(N5563), .A1(N6339), .B0(N6227));
AOI21XL inst_blk01_cellmath__39_I769 (.Y(N5944), .A0(N5898), .A1(N5901), .B0(N5706));
AOI21X1 inst_blk01_cellmath__39_I770 (.Y(N5835), .A0(N6091), .A1(N5792), .B0(N5607));
OAI2BB1X1 inst_blk01_cellmath__39_I10661 (.Y(N6020), .A0N(N5685), .A1N(N6369), .B0(N5792));
OAI21XL inst_blk01_cellmath__39_I772 (.Y(N5771), .A0(N5944), .A1(N6020), .B0(N5835));
AO21XL inst_blk01_cellmath__39_I773 (.Y(N5856), .A0(N5677), .A1(N5982), .B0(N6356));
AOI31X1 inst_blk01_cellmath__39_I10662 (.Y(N6239), .A0(N5677), .A1(N6173), .A2(N5771), .B0(N5856));
AOI21XL inst_blk01_cellmath__39_I781 (.Y(N6130), .A0(N5580), .A1(N5875), .B0(N6247));
OAI2BB1X1 inst_blk01_cellmath__39_I10663 (.Y(N6315), .A0N(N6147), .A1N(N6335), .B0(N5580));
AOI21XL inst_blk01_cellmath__39_I784 (.Y(N6015), .A0(N6325), .A1(N5758), .B0(N6138));
OAI2BB1X1 inst_blk01_cellmath__39_I10664 (.Y(N6211), .A0N(N6033), .A1N(N6222), .B0(N6325));
OA21X1 inst_blk01_cellmath__39_I790 (.Y(N6137), .A0(N6211), .A1(N6130), .B0(N6015));
OAI31X1 inst_blk01_cellmath__39_I10665 (.Y(N5704), .A0(N6211), .A1(N6315), .A2(N6239), .B0(N6137));
NOR2XL inst_blk01_cellmath__39_I822 (.Y(N6090), .A(N5921), .B(N6114));
NAND2XL inst_blk01_cellmath__39_I823 (.Y(N6279), .A(N5921), .B(N6114));
NOR2XL inst_blk01_cellmath__39_I824 (.Y(N5606), .A(N6301), .B(N5626));
NOR2XL inst_blk01_cellmath__39_I826 (.Y(N5979), .A(N5813), .B(N6001));
NAND2XL inst_blk01_cellmath__39_I827 (.Y(N6170), .A(N5813), .B(N6001));
NOR2XL inst_blk01_cellmath__39_I828 (.Y(N6355), .A(N6194), .B(N6385));
NOR2XL inst_blk01_cellmath__39_I830 (.Y(N5871), .A(N5698), .B(N5893));
NAND2X1 inst_blk01_cellmath__39_I831 (.Y(N6058), .A(N5698), .B(N5893));
NOR2X1 inst_blk01_cellmath__39_I832 (.Y(N6245), .A(N6082), .B(N6270));
NAND2X2 inst_blk01_cellmath__39_I833 (.Y(N5577), .A(N6082), .B(N6270));
NOR2XL inst_blk01_cellmath__39_I834 (.Y(N5757), .A(N5597), .B(N5785));
NAND2X2 inst_blk01_cellmath__39_I835 (.Y(N5946), .A(N5597), .B(N5785));
NOR2X2 inst_blk01_cellmath__39_I836 (.Y(N6135), .A(N5969), .B(N6162));
NOR2X1 inst_blk01_cellmath__39_I838 (.Y(N5649), .A(N6346), .B(N5668));
NAND2X4 inst_blk01_cellmath__39_I839 (.Y(N5838), .A(N6346), .B(N5668));
ADDFX1 inst_blk01_cellmath__39_I29563 (.CO(N45246), .S(N45297), .A(N45286), .B(N45242), .CI(N45270));
ADDFX1 inst_blk01_cellmath__39_I29565 (.CO(N6236), .S(N6049), .A(N45283), .B(N45249), .CI(N45297));
NOR2X1 inst_blk01_cellmath__39_I840 (.Y(N6023), .A(N5861), .B(N6049));
NAND2X2 inst_blk01_cellmath__39_I841 (.Y(N6216), .A(N5861), .B(N6049));
ADDFHXL inst_blk01_cellmath__39_I29566 (.CO(N5745), .S(N5569), .A(N45246), .B(N45239), .CI(N45259));
NOR2X1 inst_blk01_cellmath__39_I842 (.Y(N6410), .A(N5569), .B(N6236));
NAND2X4 inst_blk01_cellmath__39_I29567 (.Y(N5720), .A(N6236), .B(N5569));
NOR2X2 inst_blk01_cellmath__39_I844 (.Y(N5912), .A(N5745), .B(N5935));
NAND2X2 inst_blk01_cellmath__39_I845 (.Y(N6104), .A(N5745), .B(N5935));
NOR2X1 inst_blk01_cellmath__39_I846 (.Y(N6291), .A(N6126), .B(N6313));
NAND2X4 inst_blk01_cellmath__39_I847 (.Y(N5620), .A(N6126), .B(N6313));
NOR2X1 inst_blk01_cellmath__39_I848 (.Y(N5806), .A(N5638), .B(N5827));
NAND2X2 inst_blk01_cellmath__39_I849 (.Y(N5993), .A(N5638), .B(N5827));
NOR2X1 inst_blk01_cellmath__39_I850 (.Y(N6186), .A(N6012), .B(N6206));
NAND2X4 inst_blk01_cellmath__39_I851 (.Y(N6373), .A(N6012), .B(N6206));
NOR2X2 inst_blk01_cellmath__39_I852 (.Y(N5689), .A(N6398), .B(N5710));
NAND2X1 inst_blk01_cellmath__39_I853 (.Y(N5886), .A(N6398), .B(N5710));
NOR2X1 inst_blk01_cellmath__39_I854 (.Y(N6073), .A(N5905), .B(N6095));
NAND2X4 inst_blk01_cellmath__39_I855 (.Y(N6260), .A(N5905), .B(N6095));
NOR2X2 inst_blk01_cellmath__39_I856 (.Y(N5592), .A(N6284), .B(N5611));
NAND2X2 inst_blk01_cellmath__39_I857 (.Y(N5775), .A(N6284), .B(N5611));
NOR2X1 inst_blk01_cellmath__39_I858 (.Y(N5961), .A(N5798), .B(N5984));
NAND2X4 inst_blk01_cellmath__39_I859 (.Y(N6151), .A(N5798), .B(N5984));
NOR2X2 inst_blk01_cellmath__39_I860 (.Y(N6338), .A(N6175), .B(N6363));
NAND2X2 inst_blk01_cellmath__39_I861 (.Y(N5660), .A(N6175), .B(N6363));
NOR2X1 inst_blk01_cellmath__39_I862 (.Y(N5853), .A(N5682), .B(N5878));
NAND2X4 inst_blk01_cellmath__39_I863 (.Y(N6037), .A(N5682), .B(N5878));
NOR2X2 inst_blk01_cellmath__39_I864 (.Y(N6226), .A(N6064), .B(N6250));
NAND2X4 inst_blk01_cellmath__39_I865 (.Y(N5561), .A(N6064), .B(N6250));
NOR2XL inst_blk01_cellmath__39_I866 (.Y(N5735), .A(N5582), .B(N5763));
NAND2X4 inst_blk01_cellmath__39_I867 (.Y(N5926), .A(N5582), .B(N5763));
NOR2X2 inst_blk01_cellmath__39_I868 (.Y(N6119), .A(N5950), .B(N6142));
NAND2X1 inst_blk01_cellmath__39_I869 (.Y(N6304), .A(N5950), .B(N6142));
NOR2XL inst_blk01_cellmath__39_I870 (.Y(N5630), .A(N6330), .B(N5652));
NAND2X1 inst_blk01_cellmath__39_I871 (.Y(N5818), .A(N6330), .B(N5652));
NOR2XL inst_blk01_cellmath__39_I872 (.Y(N6005), .A(N5842), .B(N6029));
NAND2XL inst_blk01_cellmath__39_I873 (.Y(N6198), .A(N5842), .B(N6029));
NOR2XL inst_blk01_cellmath__39_I874 (.Y(N6390), .A(N6414), .B(N6219));
NAND2XL inst_blk01_cellmath__39_I875 (.Y(N5701), .A(N6414), .B(N6219));
NOR2XL inst_blk01_cellmath__39_I876 (.Y(N5897), .A(N5725), .B(N5916));
NAND2XL inst_blk01_cellmath__39_I877 (.Y(N6086), .A(N5725), .B(N5916));
NOR2XL inst_blk01_cellmath__39_I878 (.Y(N6275), .A(N6109), .B(N6296));
NAND2XL inst_blk01_cellmath__39_I879 (.Y(N5603), .A(N6109), .B(N6296));
NOR2XL inst_blk01_cellmath__39_I880 (.Y(N5788), .A(N5622), .B(N5808));
NAND2XL inst_blk01_cellmath__39_I881 (.Y(N5974), .A(N5622), .B(N5808));
NOR2XL inst_blk01_cellmath__39_I882 (.Y(N6168), .A(N5997), .B(N6191));
NAND2XL inst_blk01_cellmath__39_I883 (.Y(N6350), .A(N5997), .B(N6191));
NOR2XL inst_blk01_cellmath__39_I884 (.Y(N5673), .A(N6379), .B(N5693));
NAND2XL inst_blk01_cellmath__39_I885 (.Y(N5868), .A(N6379), .B(N5693));
NOR2XL inst_blk01_cellmath__39_I886 (.Y(N6053), .A(N5889), .B(N6078));
NAND2XL inst_blk01_cellmath__39_I887 (.Y(N6242), .A(N5889), .B(N6078));
NOR2XL inst_blk01_cellmath__39_I888 (.Y(N5573), .A(N5594), .B(N6266));
NAND2XL inst_blk01_cellmath__39_I889 (.Y(N5751), .A(N5594), .B(N6266));
NOR2XL inst_blk01_cellmath__39_I890 (.Y(N5941), .A(N5965), .B(N5779));
NAND2XL inst_blk01_cellmath__39_I891 (.Y(N6132), .A(N5965), .B(N5779));
NOR2XL inst_blk01_cellmath__39_I892 (.Y(N6319), .A(N6156), .B(N6341));
NAND2XL inst_blk01_cellmath__39_I893 (.Y(N5645), .A(N6156), .B(N6341));
NOR2XL inst_blk01_cellmath__39_I894 (.Y(N5834), .A(N6354), .B(N5663));
NAND2XL inst_blk01_cellmath__39_I895 (.Y(N6019), .A(N6354), .B(N5663));
NOR2XL inst_blk01_cellmath__39_I896 (.Y(N6213), .A(a_man[22]), .B(a_man[21]));
NAND2XL inst_blk01_cellmath__39_I897 (.Y(N6406), .A(a_man[22]), .B(a_man[21]));
AOI21X2 inst_blk01_cellmath__39_I898 (.Y(N6100), .A0(N6279), .A1(N5704), .B0(N6090));
AOI21XL inst_blk01_cellmath__39_I899 (.Y(N5989), .A0(N6170), .A1(N5606), .B0(N5979));
OAI2BB1X1 inst_blk01_cellmath__39_I10667 (.Y(N6181), .A0N(N6301), .A1N(N5626), .B0(N6170));
OAI21X4 inst_blk01_cellmath__39_I901 (.Y(N5768), .A0(N6181), .A1(N6100), .B0(N5989));
AOI21X1 inst_blk01_cellmath__39_I902 (.Y(N5658), .A0(N6058), .A1(N6355), .B0(N5871));
OAI2BB1X1 inst_blk01_cellmath__39_I10669 (.Y(N5848), .A0N(N6194), .A1N(N6385), .B0(N6058));
AOI21X2 inst_blk01_cellmath__39_I905 (.Y(N6420), .A0(N6245), .A1(N5946), .B0(N5757));
NAND2X4 inst_blk01_cellmath__39_I906 (.Y(N5731), .A(N5946), .B(N5577));
OAI21X4 inst_blk01_cellmath__39_I907 (.Y(N6195), .A0(N5731), .A1(N5658), .B0(N6420));
NOR2X4 inst_blk01_cellmath__39_I908 (.Y(N6386), .A(N5848), .B(N5731));
AOI21X4 inst_blk01_cellmath__39_I909 (.Y(N6083), .A0(N5838), .A1(N6135), .B0(N5649));
OAI2BB1X2 inst_blk01_cellmath__39_I10673 (.Y(N6271), .A0N(N5969), .A1N(N6162), .B0(N5838));
INVXL inst_blk01_cellmath__39_I911 (.Y(N6153), .A(N6216));
AOI21X4 inst_blk01_cellmath__39_I912 (.Y(N5970), .A0(N6023), .A1(N5720), .B0(N6410));
NAND2X4 inst_blk01_cellmath__39_I913 (.Y(N6164), .A(N5720), .B(N6216));
OAI21X4 inst_blk01_cellmath__39_I914 (.Y(N5747), .A0(N6164), .A1(N6083), .B0(N5970));
NOR2X4 inst_blk01_cellmath__39_I915 (.Y(N5936), .A(N6164), .B(N6271));
AOI21X4 inst_blk01_cellmath__39_I916 (.Y(N5639), .A0(N5620), .A1(N5912), .B0(N6291));
NAND2X4 inst_blk01_cellmath__39_I917 (.Y(N5830), .A(N6104), .B(N5620));
INVXL inst_blk01_cellmath__39_I918 (.Y(N6306), .A(N5993));
AOI21X4 inst_blk01_cellmath__39_I919 (.Y(N6401), .A0(N5806), .A1(N6373), .B0(N6186));
NAND2X4 inst_blk01_cellmath__39_I920 (.Y(N5712), .A(N6373), .B(N5993));
OAI21X4 inst_blk01_cellmath__39_I921 (.Y(N6176), .A0(N5712), .A1(N5639), .B0(N6401));
NOR2X4 inst_blk01_cellmath__39_I922 (.Y(N6366), .A(N5712), .B(N5830));
AOI21X4 inst_blk01_cellmath__39_I923 (.Y(N6065), .A0(N6260), .A1(N5689), .B0(N6073));
NAND2X2 inst_blk01_cellmath__39_I924 (.Y(N6251), .A(N5886), .B(N6260));
INVXL inst_blk01_cellmath__39_I925 (.Y(N5602), .A(N5775));
AOI21X4 inst_blk01_cellmath__39_I926 (.Y(N5952), .A0(N5592), .A1(N6151), .B0(N5961));
NAND2X6 inst_blk01_cellmath__39_I927 (.Y(N6143), .A(N6151), .B(N5775));
OAI21X4 inst_blk01_cellmath__39_I928 (.Y(N5726), .A0(N6143), .A1(N6065), .B0(N5952));
NOR2X6 inst_blk01_cellmath__39_I929 (.Y(N5919), .A(N6143), .B(N6251));
AOI21X4 inst_blk01_cellmath__39_I930 (.Y(N5624), .A0(N6338), .A1(N6037), .B0(N5853));
NAND2X2 inst_blk01_cellmath__39_I931 (.Y(N5809), .A(N5660), .B(N6037));
INVXL inst_blk01_cellmath__39_I932 (.Y(N5753), .A(N5561));
AOI21X2 inst_blk01_cellmath__39_I933 (.Y(N6380), .A0(N6226), .A1(N5926), .B0(N5735));
NAND2X4 inst_blk01_cellmath__39_I934 (.Y(N5694), .A(N5561), .B(N5926));
OAI21X2 inst_blk01_cellmath__39_I935 (.Y(N6158), .A0(N5694), .A1(N5624), .B0(N6380));
NOR2X4 inst_blk01_cellmath__39_I936 (.Y(N6342), .A(N5694), .B(N5809));
AOI21X2 inst_blk01_cellmath__39_I937 (.Y(N6044), .A0(N5818), .A1(N6119), .B0(N5630));
NAND2X2 inst_blk01_cellmath__39_I938 (.Y(N6232), .A(N5818), .B(N6304));
INVXL inst_blk01_cellmath__39_I939 (.Y(N6408), .A(N6198));
AOI21XL inst_blk01_cellmath__39_I940 (.Y(N5932), .A0(N5701), .A1(N6005), .B0(N6390));
NAND2X1 inst_blk01_cellmath__39_I941 (.Y(N6124), .A(N5701), .B(N6198));
OAI21X2 inst_blk01_cellmath__39_I942 (.Y(N5707), .A0(N6124), .A1(N6044), .B0(N5932));
NOR2X2 inst_blk01_cellmath__39_I943 (.Y(N5902), .A(N6124), .B(N6232));
AOI21X1 inst_blk01_cellmath__39_I944 (.Y(N5608), .A0(N5603), .A1(N5897), .B0(N6275));
NAND2XL inst_blk01_cellmath__39_I945 (.Y(N5795), .A(N5603), .B(N6086));
INVXL inst_blk01_cellmath__39_I946 (.Y(N6183), .A(N5974));
AOI21XL inst_blk01_cellmath__39_I947 (.Y(N6359), .A0(N6350), .A1(N5788), .B0(N6168));
NAND2XL inst_blk01_cellmath__39_I948 (.Y(N5679), .A(N6350), .B(N5974));
OAI21XL inst_blk01_cellmath__39_I949 (.Y(N6140), .A0(N5679), .A1(N5608), .B0(N6359));
NOR2XL inst_blk01_cellmath__39_I950 (.Y(N6327), .A(N5679), .B(N5795));
AOI21XL inst_blk01_cellmath__39_I951 (.Y(N6026), .A0(N6242), .A1(N5673), .B0(N6053));
NAND2XL inst_blk01_cellmath__39_I952 (.Y(N6217), .A(N6242), .B(N5868));
INVXL inst_blk01_cellmath__39_I953 (.Y(N5770), .A(N5573));
INVXL inst_blk01_cellmath__39_I954 (.Y(N5957), .A(N5751));
AOI21XL inst_blk01_cellmath__39_I955 (.Y(N5914), .A0(N6132), .A1(N5573), .B0(N5941));
NAND2XL inst_blk01_cellmath__39_I956 (.Y(N6107), .A(N6132), .B(N5751));
INVXL inst_blk01_cellmath__39_I957 (.Y(N5657), .A(N6026));
INVXL inst_blk01_cellmath__39_I958 (.Y(N5850), .A(N6217));
OAI21XL inst_blk01_cellmath__39_I959 (.Y(N6189), .A0(N5957), .A1(N6026), .B0(N5770));
NOR2XL inst_blk01_cellmath__39_I960 (.Y(N6376), .A(N5957), .B(N6217));
OAI21XL inst_blk01_cellmath__39_I961 (.Y(N5691), .A0(N6107), .A1(N6026), .B0(N5914));
NOR2XL inst_blk01_cellmath__39_I962 (.Y(N5887), .A(N6107), .B(N6217));
AOI21XL inst_blk01_cellmath__39_I963 (.Y(N5855), .A0(N5868), .A1(N6140), .B0(N5673));
AOI21XL inst_blk01_cellmath__39_I964 (.Y(N6228), .A0(N5850), .A1(N6140), .B0(N5657));
AOI21XL inst_blk01_cellmath__39_I965 (.Y(N5738), .A0(N6376), .A1(N6140), .B0(N6189));
AOI21XL inst_blk01_cellmath__39_I966 (.Y(N6006), .A0(N6019), .A1(N6319), .B0(N5834));
NAND2XL inst_blk01_cellmath__39_I967 (.Y(N6199), .A(N6019), .B(N5645));
INVXL inst_blk01_cellmath__39_I968 (.Y(N6387), .A(N6406));
AO21XL inst_blk01_cellmath__39_I969 (.Y(N5641), .A0(N5887), .A1(N6140), .B0(N5691));
AND2XL inst_blk01_cellmath__39_I970 (.Y(N5829), .A(N5887), .B(N6327));
INVX1 inst_blk01_cellmath__39_I971 (.Y(N6014), .A(N5768));
AOI21X4 inst_blk01_cellmath__39_I972 (.Y(N6102), .A0(N6386), .A1(N5768), .B0(N6195));
AOI21X4 inst_blk01_cellmath__39_I973 (.Y(N5617), .A0(N5936), .A1(N6195), .B0(N5747));
NAND2X4 inst_blk01_cellmath__39_I974 (.Y(N5804), .A(N5936), .B(N6386));
AOI21X4 inst_blk01_cellmath__39_I975 (.Y(N5991), .A0(N6366), .A1(N5747), .B0(N6176));
NAND2X4 inst_blk01_cellmath__39_I976 (.Y(N6184), .A(N6366), .B(N5936));
AOI21X4 inst_blk01_cellmath__39_I977 (.Y(N6371), .A0(N5919), .A1(N6176), .B0(N5726));
NAND2X4 inst_blk01_cellmath__39_I978 (.Y(N5688), .A(N6366), .B(N5919));
AOI21X4 inst_blk01_cellmath__39_I979 (.Y(N5884), .A0(N6342), .A1(N5726), .B0(N6158));
NAND2X4 inst_blk01_cellmath__39_I980 (.Y(N6071), .A(N6342), .B(N5919));
AOI21X2 inst_blk01_cellmath__39_I981 (.Y(N6258), .A0(N5902), .A1(N6158), .B0(N5707));
NAND2X2 inst_blk01_cellmath__39_I982 (.Y(N5590), .A(N5902), .B(N6342));
AOI21X1 inst_blk01_cellmath__39_I983 (.Y(N5773), .A0(N5829), .A1(N5707), .B0(N5641));
NAND2X2 inst_blk01_cellmath__39_I984 (.Y(N5959), .A(N5829), .B(N5902));
INVXL inst_blk01_cellmath__39_I985 (.Y(N6208), .A(N6014));
INVX1 inst_blk01_cellmath__39_I986 (.Y(N6400), .A(N6102));
OAI21X4 inst_blk01_cellmath__39_I987 (.Y(N6035), .A0(N5804), .A1(N6014), .B0(N5617));
OAI21X4 inst_blk01_cellmath__39_I988 (.Y(N5559), .A0(N6102), .A1(N6184), .B0(N5991));
OAI21X1 inst_blk01_cellmath__39_I989 (.Y(N5924), .A0(N5688), .A1(N5617), .B0(N6371));
NOR2X1 inst_blk01_cellmath__39_I990 (.Y(N6116), .A(N5688), .B(N5804));
OAI21X2 inst_blk01_cellmath__39_I991 (.Y(N6302), .A0(N6071), .A1(N5991), .B0(N5884));
NOR2X1 inst_blk01_cellmath__39_I992 (.Y(N5628), .A(N6071), .B(N6184));
OAI21X4 inst_blk01_cellmath__39_I993 (.Y(N5816), .A0(N5590), .A1(N6371), .B0(N6258));
NOR2X2 inst_blk01_cellmath__39_I994 (.Y(N6003), .A(N5688), .B(N5590));
OAI21X4 inst_blk01_cellmath__39_I995 (.Y(N6196), .A0(N5959), .A1(N5884), .B0(N5773));
NOR2X2 inst_blk01_cellmath__39_I996 (.Y(N6389), .A(N5959), .B(N6071));
INVXL inst_blk01_cellmath__39_I999 (.Y(N6097), .A(N6035));
INVXL inst_blk01_cellmath__39_I1000 (.Y(N6286), .A(N5559));
AOI21X2 inst_blk01_cellmath__39_I1001 (.Y(N6349), .A0(N6116), .A1(N6208), .B0(N5924));
NOR2XL inst_blk01_cellmath__39_I1009 (.Y(N5928), .A(N6153), .B(N6083));
NOR2XL inst_blk01_cellmath__39_I1010 (.Y(N5844), .A(N5928), .B(N6023));
NOR2XL inst_blk01_cellmath__39_I1011 (.Y(N6393), .A(N6306), .B(N5639));
NOR2XL inst_blk01_cellmath__39_I1012 (.Y(N6111), .A(N6393), .B(N5806));
NOR2XL inst_blk01_cellmath__39_I1013 (.Y(N6394), .A(N5602), .B(N6065));
NOR2XL inst_blk01_cellmath__39_I1014 (.Y(N6382), .A(N5592), .B(N6394));
NOR2X1 inst_blk01_cellmath__39_I1015 (.Y(N5977), .A(N5753), .B(N5624));
NOR2XL inst_blk01_cellmath__39_I1016 (.Y(N5781), .A(N5977), .B(N6226));
NOR2XL inst_blk01_cellmath__39_I1017 (.Y(N5576), .A(N6408), .B(N6044));
NOR2XL inst_blk01_cellmath__39_I1018 (.Y(N6046), .A(N5576), .B(N6005));
NOR2XL inst_blk01_cellmath__39_I1019 (.Y(N6022), .A(N6183), .B(N5608));
NOR2XL inst_blk01_cellmath__39_I1020 (.Y(N6311), .A(N6022), .B(N5788));
INVXL inst_blk01_cellmath__39_I1021 (.Y(N5825), .A(N6140));
NOR2XL inst_blk01_cellmath__39_I1022 (.Y(N5619), .A(N6387), .B(N6006));
NOR2XL inst_blk01_cellmath__39_I1023 (.Y(N6358), .A(N5619), .B(N6213));
OR2XL inst_blk01_cellmath__39_I1024 (.Y(N5681), .A(N6387), .B(N6199));
NAND2BXL inst_blk01_cellmath__39_I1035 (.Y(N5564), .AN(N6410), .B(N5720));
NAND2BXL inst_blk01_cellmath__39_I1036 (.Y(N6412), .AN(N5912), .B(N6104));
NAND2BXL inst_blk01_cellmath__39_I1037 (.Y(N6106), .AN(N6291), .B(N5620));
NAND2BXL inst_blk01_cellmath__39_I1038 (.Y(N6353), .AN(N5806), .B(N5993));
NAND2BXL inst_blk01_cellmath__39_I1039 (.Y(N5836), .AN(N6186), .B(N6373));
NAND2BXL inst_blk01_cellmath__39_I1040 (.Y(N6075), .AN(N5689), .B(N5886));
NAND2BXL inst_blk01_cellmath__39_I1041 (.Y(N5777), .AN(N6073), .B(N6260));
NAND2BXL inst_blk01_cellmath__39_I1042 (.Y(N5772), .AN(N5592), .B(N5775));
NAND2BXL inst_blk01_cellmath__39_I1043 (.Y(N6118), .AN(N5961), .B(N6151));
NAND2BXL inst_blk01_cellmath__39_I1044 (.Y(N5737), .AN(N6338), .B(N5660));
NAND2BXL inst_blk01_cellmath__39_I1045 (.Y(N6307), .AN(N5853), .B(N6037));
NAND2BXL inst_blk01_cellmath__39_I1046 (.Y(N6052), .AN(N6226), .B(N5561));
NAND2BXL inst_blk01_cellmath__39_I1047 (.Y(N6404), .AN(N5735), .B(N5926));
NAND2BXL inst_blk01_cellmath__39_I1048 (.Y(N6277), .AN(N6119), .B(N6304));
NAND2BXL inst_blk01_cellmath__39_I1049 (.Y(N5975), .AN(N5630), .B(N5818));
NAND2BXL inst_blk01_cellmath__39_I1050 (.Y(N6334), .AN(N6005), .B(N6198));
NAND2BXL inst_blk01_cellmath__39_I1051 (.Y(N5814), .AN(N6390), .B(N5701));
NAND2BXL inst_blk01_cellmath__39_I1053 (.Y(N5647), .AN(N6275), .B(N5603));
NAND2BXL inst_blk01_cellmath__39_I1054 (.Y(N5746), .AN(N5788), .B(N5974));
NAND2BXL inst_blk01_cellmath__39_I1055 (.Y(N6094), .AN(N6168), .B(N6350));
NAND2BXL inst_blk01_cellmath__39_I1056 (.Y(N5583), .AN(N5673), .B(N5868));
NAND2BXL inst_blk01_cellmath__39_I1057 (.Y(N5917), .AN(N6053), .B(N6242));
NAND2BXL inst_blk01_cellmath__39_I1058 (.Y(N6265), .AN(N5573), .B(N5751));
NAND2BXL inst_blk01_cellmath__39_I1059 (.Y(N5741), .AN(N5941), .B(N6132));
NAND2BXL inst_blk01_cellmath__39_I1061 (.Y(N5851), .AN(N5834), .B(N6019));
NAND2BXL inst_blk01_cellmath__39_I1062 (.Y(N5678), .AN(N6213), .B(N6406));
XNOR2X1 inst_blk01_cellmath__39_I1068 (.Y(N624), .A(N6097), .B(N6412));
XNOR2X1 inst_blk01_cellmath__39_I1069 (.Y(N628), .A(N6075), .B(N6286));
XNOR2X1 inst_blk01_cellmath__39_I1070 (.Y(N632), .A(N5737), .B(N6349));
AOI21X2 inst_cellmath__48_I29633 (.Y(N5865), .A0(N5628), .A1(N6400), .B0(N6302));
XNOR2X1 inst_blk01_cellmath__39_I1071 (.Y(N636), .A(N6277), .B(N5865));
XOR2XL inst_blk01_cellmath__39_I1093 (.Y(N5643), .A(N5564), .B(N5844));
OAI21XL inst_blk01_cellmath__39_I1094 (.Y(N6040), .A0(N6153), .A1(N6271), .B0(N5844));
XNOR2X1 inst_blk01_cellmath__39_I1095 (.Y(N5832), .A(N5564), .B(N6040));
MXI2XL inst_blk01_cellmath__39_I1096 (.Y(N623), .A(N5643), .B(N5832), .S0(N6400));
XNOR2X1 inst_blk01_cellmath__39_I1097 (.Y(N6403), .A(N6106), .B(N6104));
XNOR2X1 inst_blk01_cellmath__39_I1098 (.Y(N6210), .A(N5912), .B(N6106));
MXI2XL inst_blk01_cellmath__39_I1099 (.Y(N625), .A(N6403), .B(N6210), .S0(N6097));
XOR2XL inst_blk01_cellmath__39_I1100 (.Y(N5909), .A(N5639), .B(N6353));
NAND2XL inst_blk01_cellmath__39_I1101 (.Y(N5978), .A(N5830), .B(N5639));
XNOR2X1 inst_blk01_cellmath__39_I1102 (.Y(N6099), .A(N6353), .B(N5978));
MXI2XL inst_blk01_cellmath__39_I1103 (.Y(N626), .A(N6099), .B(N5909), .S0(N6097));
XOR2XL inst_blk01_cellmath__39_I1104 (.Y(N5614), .A(N5836), .B(N6111));
OAI21XL inst_blk01_cellmath__39_I1105 (.Y(N6321), .A0(N6306), .A1(N5830), .B0(N6111));
INVXL xnor2_A_I30573 (.Y(N45756), .A(N5836));
MXI2XL xnor2_A_I30574 (.Y(N5801), .A(N5836), .B(N45756), .S0(N6321));
MXI2XL inst_blk01_cellmath__39_I1107 (.Y(N627), .A(N5801), .B(N5614), .S0(N6097));
XNOR2X1 inst_blk01_cellmath__39_I1108 (.Y(N6368), .A(N5886), .B(N5777));
XNOR2X1 inst_blk01_cellmath__39_I1109 (.Y(N6179), .A(N5689), .B(N5777));
MXI2XL inst_blk01_cellmath__39_I10403 (.Y(N23218), .A(N6368), .B(N6179), .S0(N6286));
XOR2XL inst_blk01_cellmath__39_I1111 (.Y(N5881), .A(N6065), .B(N5772));
NAND2XL inst_blk01_cellmath__39_I1112 (.Y(N6257), .A(N6251), .B(N6065));
XNOR2X1 inst_blk01_cellmath__39_I1113 (.Y(N6068), .A(N5772), .B(N6257));
MXI2XL inst_blk01_cellmath__39_I1114 (.Y(N630), .A(N6068), .B(N5881), .S0(N6286));
XOR2XL inst_blk01_cellmath__39_I1115 (.Y(N5587), .A(N6382), .B(N6118));
OAI21XL inst_blk01_cellmath__39_I1116 (.Y(N5733), .A0(N5602), .A1(N6251), .B0(N6382));
XNOR2XL inst_blk01_cellmath__39_I1117 (.Y(N5766), .A(N6118), .B(N5733));
MXI2X1 inst_blk01_cellmath__39_I1118 (.Y(N631), .A(N5766), .B(N5587), .S0(N6286));
XNOR2X1 inst_blk01_cellmath__39_I1119 (.Y(N6333), .A(N6307), .B(N5660));
XNOR2X1 inst_blk01_cellmath__39_I1120 (.Y(N6146), .A(N6307), .B(N6338));
MXI2XL inst_blk01_cellmath__39_I1121 (.Y(N633), .A(N6333), .B(N6146), .S0(N6349));
XOR2XL inst_blk01_cellmath__39_I1122 (.Y(N5846), .A(N6052), .B(N5624));
NAND2XL inst_blk01_cellmath__39_I1123 (.Y(N5672), .A(N5809), .B(N5624));
XNOR2X1 inst_blk01_cellmath__39_I1124 (.Y(N6032), .A(N6052), .B(N5672));
MXI2XL inst_blk01_cellmath__39_I1125 (.Y(N634), .A(N6032), .B(N5846), .S0(N6349));
XOR2XL inst_blk01_cellmath__39_I1126 (.Y(N6418), .A(N6404), .B(N5781));
OAI21XL inst_blk01_cellmath__39_I1127 (.Y(N6018), .A0(N5753), .A1(N5809), .B0(N5781));
XNOR2XL inst_blk01_cellmath__39_I1128 (.Y(N5729), .A(N6404), .B(N6018));
MXI2XL inst_blk01_cellmath__39_I1129 (.Y(N635), .A(N5729), .B(N6418), .S0(N6349));
XNOR2X1 inst_blk01_cellmath__39_I1130 (.Y(N6299), .A(N5975), .B(N6304));
XNOR2X1 inst_blk01_cellmath__39_I1131 (.Y(N6112), .A(N5975), .B(N6119));
MXI2XL inst_blk01_cellmath__39_I1132 (.Y(N637), .A(N6299), .B(N6112), .S0(N5865));
NAND2XL inst_blk01_cellmath__39_I1134 (.Y(N5955), .A(N6232), .B(N6044));
OAI21XL inst_blk01_cellmath__39_I1138 (.Y(N6300), .A0(N6408), .A1(N6232), .B0(N6046));
XOR2XL inst_blk01_cellmath__39_I1144 (.Y(N5784), .A(N5746), .B(N5608));
NAND2XL inst_blk01_cellmath__39_I1145 (.Y(N6235), .A(N5795), .B(N5608));
XNOR2X1 inst_blk01_cellmath__39_I1146 (.Y(N5968), .A(N5746), .B(N6235));
AOI21X4 inst_cellmath__48_I29637 (.Y(N6240), .A0(N6003), .A1(N6035), .B0(N5816));
MXI2XL inst_blk01_cellmath__39_I1147 (.Y(N642), .A(N5968), .B(N5784), .S0(N6240));
XOR2XL inst_blk01_cellmath__39_I1148 (.Y(N6345), .A(N6094), .B(N6311));
OAI21XL inst_blk01_cellmath__39_I1149 (.Y(N5711), .A0(N6183), .A1(N5795), .B0(N6311));
XNOR2X1 inst_blk01_cellmath__39_I1150 (.Y(N5666), .A(N6094), .B(N5711));
MXI2X1 inst_blk01_cellmath__39_I1151 (.Y(N643), .A(N5666), .B(N6345), .S0(N6240));
XOR2XL inst_blk01_cellmath__39_I1152 (.Y(N6048), .A(N5583), .B(N5825));
NAND2BXL inst_blk01_cellmath__39_I1153 (.Y(N6063), .AN(N6327), .B(N5825));
XNOR2X1 inst_blk01_cellmath__39_I1154 (.Y(N6234), .A(N5583), .B(N6063));
MXI2X1 inst_blk01_cellmath__39_I1155 (.Y(N644), .A(N6234), .B(N6048), .S0(N6240));
XOR2XL inst_blk01_cellmath__39_I1156 (.Y(N5744), .A(N5917), .B(N5855));
OAI2BB1X1 inst_blk01_cellmath__39_I1157 (.Y(N6415), .A0N(N5868), .A1N(N6327), .B0(N5855));
XNOR2X1 inst_blk01_cellmath__39_I1158 (.Y(N5934), .A(N5917), .B(N6415));
MXI2XL inst_blk01_cellmath__39_I1159 (.Y(N645), .A(N5934), .B(N5744), .S0(N6240));
OAI2BB1X1 inst_blk01_cellmath__39_I1161 (.Y(N5890), .A0N(N5850), .A1N(N6327), .B0(N6228));
OAI2BB1X1 inst_blk01_cellmath__39_I1165 (.Y(N6230), .A0N(N6376), .A1N(N6327), .B0(N5738));
XOR2XL inst_blk01_cellmath__39_I1171 (.Y(N6283), .A(N5678), .B(N6006));
NAND2XL inst_blk01_cellmath__39_I1172 (.Y(N6172), .A(N6199), .B(N6006));
XNOR2X1 inst_blk01_cellmath__39_I1173 (.Y(N5610), .A(N5678), .B(N6172));
AOI21X4 inst_cellmath__48_I29461 (.Y(N5750), .A0(N6389), .A1(N5559), .B0(N6196));
MXI2X1 inst_blk01_cellmath__39_I1174 (.Y(N650), .A(N5610), .B(N6283), .S0(N5750));
OA21XL inst_blk01_cellmath__39_I1175 (.Y(N652), .A0(N5681), .A1(N5750), .B0(N6358));
INVX1 inst_blk01_cellmath__39_I1176 (.Y(N651), .A(N652));
INVXL inst_cellmath__42_0_I1179 (.Y(N7287), .A(a_exp[2]));
INVXL inst_cellmath__42_0_I1180 (.Y(N7293), .A(a_exp[3]));
INVXL inst_cellmath__42_0_I1181 (.Y(N7264), .A(a_exp[4]));
INVXL inst_cellmath__42_0_I1183 (.Y(N7268), .A(a_exp[6]));
INVXL inst_cellmath__48_I29650 (.Y(N7280), .A(a_exp[1]));
OAI21XL inst_cellmath__42_0_I1184 (.Y(N7284), .A0(N7287), .A1(N7280), .B0(N7293));
INVXL inst_cellmath__48_I29441 (.Y(N7289), .A(a_exp[5]));
NAND3XL inst_cellmath__42_0_I1185 (.Y(N7281), .A(N7268), .B(N7289), .C(N7264));
INVXL inst_cellmath__42_0_I1186 (.Y(N7267), .A(a_exp[7]));
NAND2XL inst_cellmath__42_0_I1187 (.Y(N7270), .A(N7289), .B(N7264));
NOR2XL inst_cellmath__42_0_I1188 (.Y(N7271), .A(N7284), .B(N7270));
NOR2XL node_cs_const1_cs_A_I30575 (.Y(N45763), .A(N7287), .B(N7280));
XNOR2X1 node_cs_const1_cs_A_I30576 (.Y(inst_cellmath__42[3]), .A(N7293), .B(N45763));
XOR2XL inst_cellmath__42_0_I1196 (.Y(inst_cellmath__42[6]), .A(N7271), .B(N7268));
NOR2XL inst_cellmath__42_0_I1197 (.Y(N7291), .A(N7281), .B(N7284));
XNOR2X1 inst_cellmath__42_0_I1198 (.Y(inst_cellmath__42[7]), .A(N7267), .B(N7291));
MXI2XL inst_cellmath__48_I1209 (.Y(N7360), .A(N624), .B(N623), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1210 (.Y(N7418), .A(N625), .B(N624), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1211 (.Y(N7472), .A(N626), .B(N625), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1212 (.Y(N7529), .A(N627), .B(N626), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1213 (.Y(N7329), .A(N628), .B(N627), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1214 (.Y(N7385), .A(N23218), .B(N628), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1215 (.Y(N7441), .A(N630), .B(N23218), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1216 (.Y(N7495), .A(N631), .B(N630), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1217 (.Y(N7551), .A(N632), .B(N631), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1218 (.Y(N7351), .A(N633), .B(N632), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1219 (.Y(N7408), .A(N634), .B(N633), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1220 (.Y(N7463), .A(N635), .B(N634), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1221 (.Y(N7519), .A(N636), .B(N635), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1222 (.Y(N7321), .A(N637), .B(N636), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I29640 (.Y(N45460), .A(N6334), .B(N5955));
XOR2XL inst_cellmath__48_I29639 (.Y(N45451), .A(N6334), .B(N6044));
MXI2XL inst_cellmath__48_I29641 (.Y(N638), .A(N45460), .B(N45451), .S0(N5865));
MXI2XL inst_cellmath__48_I1223 (.Y(N7373), .A(N638), .B(N637), .S0(a_exp[0]));
NOR2BX1 inst_cellmath__48_I29727 (.Y(N45456), .AN(N6086), .B(N5897));
INVXL inst_cellmath__48_I29636 (.Y(N45454), .A(N45456));
MXI2XL inst_cellmath__48_I29638 (.Y(N640), .A(N45454), .B(N45456), .S0(N6240));
XNOR2X1 inst_cellmath__48_I29643 (.Y(N45446), .A(N5814), .B(N6300));
XOR2XL inst_cellmath__48_I29642 (.Y(N45439), .A(N5814), .B(N6046));
MXI2X1 inst_cellmath__48_I29644 (.Y(N639), .A(N45446), .B(N45439), .S0(N5865));
MXI2XL inst_cellmath__48_I1225 (.Y(N7486), .A(N640), .B(N639), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I29645 (.Y(N45464), .A(N5647), .B(N6086));
XNOR2X1 inst_cellmath__48_I29646 (.Y(N45473), .A(N5647), .B(N5897));
MXI2XL inst_cellmath__48_I29647 (.Y(N641), .A(N45464), .B(N45473), .S0(N6240));
MXI2XL inst_cellmath__48_I1227 (.Y(N7344), .A(N642), .B(N641), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1228 (.Y(N7401), .A(N643), .B(N642), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1229 (.Y(N7454), .A(N644), .B(N643), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1230 (.Y(N7508), .A(N645), .B(N644), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I29469 (.Y(N45061), .A(N6265), .B(N5890));
XOR2XL inst_cellmath__48_I29468 (.Y(N45051), .A(N6265), .B(N6228));
MXI2XL inst_cellmath__48_I29470 (.Y(N646), .A(N45061), .B(N45051), .S0(N6240));
MXI2X1 inst_cellmath__48_I1231 (.Y(N7565), .A(N646), .B(N645), .S0(a_exp[0]));
NAND2BXL inst_cellmath__48_I29462 (.Y(N45027), .AN(N6319), .B(N5645));
XNOR2X1 inst_cellmath__48_I29467 (.Y(N648), .A(N45027), .B(N5750));
XNOR2X1 inst_cellmath__48_I29472 (.Y(N45046), .A(N5741), .B(N6230));
XOR2XL inst_cellmath__48_I29471 (.Y(N45032), .A(N5741), .B(N5738));
MXI2XL inst_cellmath__48_I29473 (.Y(N647), .A(N45046), .B(N45032), .S0(N6240));
MXI2XL inst_cellmath__48_I1233 (.Y(N7424), .A(N648), .B(N647), .S0(a_exp[0]));
XNOR2X1 inst_cellmath__48_I29474 (.Y(N45067), .A(N5851), .B(N5645));
XNOR2X1 inst_cellmath__48_I29475 (.Y(N45025), .A(N5851), .B(N6319));
MXI2XL inst_cellmath__48_I29481 (.Y(N649), .A(N45067), .B(N45025), .S0(N5750));
MXI2XL inst_cellmath__48_I1235 (.Y(N7533), .A(N650), .B(N649), .S0(a_exp[0]));
MXI2X1 inst_cellmath__48_I1236 (.Y(N7333), .A(N651), .B(N650), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I1237 (.Y(N7391), .A(N652), .B(N651), .S0(a_exp[0]));
NAND2XL inst_cellmath__48_I1238 (.Y(N7447), .A(N652), .B(a_exp[0]));
INVXL inst_cellmath__48_I29463 (.Y(N45023), .A(N5750));
NAND2XL inst_cellmath__48_I29464 (.Y(N45020), .A(N45027), .B(N5750));
NAND2BXL inst_cellmath__48_I29729 (.Y(N45072), .AN(N45027), .B(N45023));
INVXL inst_cellmath__48_I29477 (.Y(N45068), .A(N5750));
NOR2BX1 inst_cellmath__48_I29730 (.Y(N45033), .AN(N45025), .B(N45068));
INVXL inst_cellmath__48_I29479 (.Y(N45040), .A(N45067));
NOR2XL inst_cellmath__48_I29480 (.Y(N45050), .A(N45040), .B(N5750));
MXI2XL inst_cellmath__48_I29648 (.Y(N7432), .A(N639), .B(N638), .S0(a_exp[0]));
MXI2XL inst_cellmath__48_I29649 (.Y(N7543), .A(N641), .B(N640), .S0(a_exp[0]));
CLKINVX12 inst_cellmath__48_I29651 (.Y(inst_cellmath__42[1]), .A(N7280));
MXI2XL inst_cellmath__48_I29652 (.Y(N7475), .A(N7432), .B(N7543), .S0(a_exp[1]));
INVX1 inst_cellmath__48_I29484 (.Y(N45071), .A(a_exp[0]));
INVXL inst_cellmath__48_I29485 (.Y(N45019), .A(N45061));
INVXL inst_cellmath__48_I29486 (.Y(N45064), .A(N45051));
MXI2XL inst_cellmath__48_I29487 (.Y(N45045), .A(N45019), .B(N45064), .S0(N6240));
NOR2XL inst_cellmath__48_I29488 (.Y(N45070), .A(N45071), .B(N45045));
INVXL inst_cellmath__48_I29489 (.Y(N45016), .A(N45046));
INVXL inst_cellmath__48_I29490 (.Y(N45043), .A(N45032));
MXI2XL inst_cellmath__48_I29491 (.Y(N45065), .A(N45016), .B(N45043), .S0(N6240));
NOR2X1 inst_cellmath__48_I29492 (.Y(N45031), .A(a_exp[0]), .B(N45065));
MXI2XL inst_cellmath__48_I29493 (.Y(N7365), .A(N647), .B(N646), .S0(a_exp[0]));
AOI21X1 inst_cellmath__48_I29494 (.Y(N45036), .A0(N45072), .A1(N45020), .B0(N45071));
NOR3X1 inst_cellmath__48_I29495 (.Y(N45052), .A(a_exp[0]), .B(N45050), .C(N45033));
MXI2XL inst_cellmath__48_I29496 (.Y(N7478), .A(N649), .B(N648), .S0(a_exp[0]));
NOR3BXL inst_cellmath__48_I29735 (.Y(N45055), .AN(inst_cellmath__42[1]), .B(N45052), .C(N45036));
NOR3X1 inst_cellmath__48_I29499 (.Y(N45015), .A(inst_cellmath__42[1]), .B(N45070), .C(N45031));
NOR2XL inst_cellmath__48_I29500 (.Y(N7411), .A(N45015), .B(N45055));
MXI2XL inst_cellmath__48_I1246 (.Y(N7407), .A(N7360), .B(N7472), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1247 (.Y(N7462), .A(N7418), .B(N7529), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1248 (.Y(N7516), .A(N7472), .B(N7329), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1249 (.Y(N7318), .A(N7529), .B(N7385), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1250 (.Y(N7372), .A(N7329), .B(N7441), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1251 (.Y(N7431), .A(N7385), .B(N7495), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1252 (.Y(N7484), .A(N7441), .B(N7551), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1253 (.Y(N7541), .A(N7495), .B(N7351), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1254 (.Y(N7341), .A(N7551), .B(N7408), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1255 (.Y(N7398), .A(N7351), .B(N7463), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1256 (.Y(N7453), .A(N7408), .B(N7519), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1257 (.Y(N7507), .A(N7463), .B(N7321), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1258 (.Y(N7563), .A(N7519), .B(N7373), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1259 (.Y(N7363), .A(N7321), .B(N7432), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1260 (.Y(N7421), .A(N7373), .B(N7486), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1262 (.Y(N7532), .A(N7486), .B(N7344), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1263 (.Y(N7332), .A(N7543), .B(N7401), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1264 (.Y(N7388), .A(N7344), .B(N7454), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1265 (.Y(N7444), .A(N7401), .B(N7508), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1266 (.Y(N7499), .A(N7454), .B(N7565), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1267 (.Y(N7554), .A(N7508), .B(N7365), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1268 (.Y(N7354), .A(N7565), .B(N7424), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1270 (.Y(N7467), .A(N7424), .B(N7533), .S0(inst_cellmath__42[1]));
MXI2X1 inst_cellmath__48_I1271 (.Y(N7522), .A(N7478), .B(N7333), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1272 (.Y(N7325), .A(N7533), .B(N7391), .S0(inst_cellmath__42[1]));
MXI2XL inst_cellmath__48_I1273 (.Y(N7378), .A(N7333), .B(N7447), .S0(inst_cellmath__42[1]));
NOR2XL inst_cellmath__48_I1274 (.Y(N7437), .A(inst_cellmath__42[1]), .B(N7391));
NOR2XL inst_cellmath__48_I1275 (.Y(N7547), .A(inst_cellmath__42[1]), .B(N7447));
CLKMX2X6 inst_cellmath__48_I10677 (.Y(N7468), .A(N7280), .B(inst_cellmath__42[1]), .S0(N7287));
MXI2XL inst_cellmath__48_I1284 (.Y(N7506), .A(N7372), .B(N7407), .S0(N7468));
MXI2XL inst_cellmath__48_I1285 (.Y(N7562), .A(N7431), .B(N7462), .S0(N7468));
MXI2XL inst_cellmath__48_I1286 (.Y(N7362), .A(N7484), .B(N7516), .S0(N7468));
MXI2XL inst_cellmath__48_I1287 (.Y(N7419), .A(N7541), .B(N7318), .S0(N7468));
MXI2XL inst_cellmath__48_I1288 (.Y(N7473), .A(N7341), .B(N7372), .S0(N7468));
MXI2XL inst_cellmath__48_I1289 (.Y(N7531), .A(N7398), .B(N7431), .S0(N7468));
MXI2XL inst_cellmath__48_I1290 (.Y(N7331), .A(N7453), .B(N7484), .S0(N7468));
MXI2XL inst_cellmath__48_I1291 (.Y(N7387), .A(N7507), .B(N7541), .S0(N7468));
MXI2X1 inst_cellmath__48_I1292 (.Y(N7443), .A(N7563), .B(N7341), .S0(N7468));
MXI2X1 inst_cellmath__48_I1293 (.Y(N7496), .A(N7363), .B(N7398), .S0(N7468));
MXI2X1 inst_cellmath__48_I1294 (.Y(N7552), .A(N7421), .B(N7453), .S0(N7468));
MXI2XL inst_cellmath__48_I1295 (.Y(N7353), .A(N7475), .B(N7507), .S0(N7468));
MXI2XL inst_cellmath__48_I1296 (.Y(N7410), .A(N7532), .B(N7563), .S0(N7468));
MXI2XL inst_cellmath__48_I1297 (.Y(N7466), .A(N7332), .B(N7363), .S0(N7468));
MXI2X1 inst_cellmath__48_I1298 (.Y(N7521), .A(N7388), .B(N7421), .S0(N7468));
MXI2XL inst_cellmath__48_I1299 (.Y(N7322), .A(N7444), .B(N7475), .S0(N7468));
MXI2X1 inst_cellmath__48_I1300 (.Y(N7376), .A(N7499), .B(N7532), .S0(N7468));
MXI2X1 inst_cellmath__48_I1301 (.Y(N7436), .A(N7554), .B(N7332), .S0(N7468));
MXI2X1 inst_cellmath__48_I1302 (.Y(N7489), .A(N7354), .B(N7388), .S0(N7468));
MXI2XL inst_cellmath__48_I1303 (.Y(N7546), .A(N7411), .B(N7444), .S0(N7468));
MXI2XL inst_cellmath__48_I1304 (.Y(N7346), .A(N7467), .B(N7499), .S0(N7468));
MXI2XL inst_cellmath__48_I1305 (.Y(N7402), .A(N7522), .B(N7554), .S0(N7468));
MXI2XL inst_cellmath__48_I1306 (.Y(N7457), .A(N7325), .B(N7354), .S0(N7468));
MXI2X1 inst_cellmath__48_I1307 (.Y(N7512), .A(N7378), .B(N7411), .S0(N7468));
MXI2X1 inst_cellmath__48_I1308 (.Y(N7568), .A(N7437), .B(N7467), .S0(N7468));
MXI2XL inst_cellmath__48_I1309 (.Y(N7368), .A(N7547), .B(N7522), .S0(N7468));
NAND2XL inst_cellmath__48_I1310 (.Y(N7426), .A(N7468), .B(N7325));
NAND2XL inst_cellmath__48_I1311 (.Y(N7536), .A(N7468), .B(N7378));
NAND2XL inst_cellmath__48_I1312 (.Y(N7394), .A(N7437), .B(N7468));
NAND2XL inst_cellmath__48_I1313 (.Y(N7503), .A(N7547), .B(N7468));
MXI2XL inst_cellmath__48_I1324 (.Y(N7464), .A(N7506), .B(N7443), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1325 (.Y(N7518), .A(N7562), .B(N7496), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1326 (.Y(N7320), .A(N7362), .B(N7552), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1327 (.Y(N7375), .A(N7419), .B(N7353), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1328 (.Y(N7434), .A(N7473), .B(N7410), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1329 (.Y(N7487), .A(N7531), .B(N7466), .S0(inst_cellmath__42[3]));
MXI2X1 inst_cellmath__48_I1330 (.Y(N7544), .A(N7331), .B(N7521), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1331 (.Y(N7343), .A(N7387), .B(N7322), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1332 (.Y(N7400), .A(N7443), .B(N7376), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1333 (.Y(N7456), .A(N7496), .B(N7436), .S0(inst_cellmath__42[3]));
MXI2X1 inst_cellmath__48_I1334 (.Y(N7510), .A(N7552), .B(N7489), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1335 (.Y(N7566), .A(N7353), .B(N7546), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1336 (.Y(N7366), .A(N7410), .B(N7346), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1337 (.Y(N7423), .A(N7466), .B(N7402), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1338 (.Y(N7477), .A(N7521), .B(N7457), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1339 (.Y(N7535), .A(N7322), .B(N7512), .S0(inst_cellmath__42[3]));
MXI2X1 inst_cellmath__48_I1340 (.Y(N7335), .A(N7376), .B(N7568), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1341 (.Y(N7392), .A(N7436), .B(N7368), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1342 (.Y(N7448), .A(N7489), .B(N7426), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1343 (.Y(N7501), .A(N7546), .B(N7536), .S0(inst_cellmath__42[3]));
MXI2XL inst_cellmath__48_I1344 (.Y(N7557), .A(N7346), .B(N7394), .S0(inst_cellmath__42[3]));
MXI2X1 inst_cellmath__48_I1345 (.Y(N7357), .A(N7402), .B(N7503), .S0(inst_cellmath__42[3]));
NOR2X1 inst_cellmath__48_I1346 (.Y(N7414), .A(inst_cellmath__42[3]), .B(N7457));
NOR2XL inst_cellmath__48_I1348 (.Y(N7381), .A(N7568), .B(inst_cellmath__42[3]));
NOR2XL inst_cellmath__48_I1349 (.Y(N7492), .A(inst_cellmath__42[3]), .B(N7368));
NOR2XL inst_cellmath__48_I1350 (.Y(N7349), .A(N7426), .B(inst_cellmath__42[3]));
NOR2XL inst_cellmath__48_I1351 (.Y(N7460), .A(N7536), .B(inst_cellmath__42[3]));
NOR2X1 inst_cellmath__48_I1352 (.Y(N7570), .A(inst_cellmath__42[3]), .B(N7394));
NOR2XL inst_cellmath__48_I1353 (.Y(N7428), .A(N7503), .B(inst_cellmath__42[3]));
NOR2XL inst_cellmath__48_I29442 (.Y(N44974), .A(a_exp[4]), .B(N7284));
XNOR2X1 inst_cellmath__48_I30072 (.Y(N44981), .A(N44974), .B(N7289));
XOR2X4 inst_cellmath__48_I29448 (.Y(N7395), .A(N7264), .B(N7284));
MXI2XL inst_cellmath__48_I29654 (.Y(N45504), .A(N7460), .B(N7566), .S0(N7395));
XOR2X4 inst_cellmath__48_I29655 (.Y(inst_cellmath__42[5]), .A(N7289), .B(N44974));
NOR2XL inst_cellmath__48_I29656 (.Y(N45494), .A(inst_cellmath__42[5]), .B(N45504));
NOR2X2 inst_cellmath__48_I29447 (.Y(N7525), .A(inst_cellmath__42[3]), .B(N7512));
NAND3X4 inst_cellmath__48_I29451 (.Y(N7812), .A(N44981), .B(N7395), .C(N7525));
INVX3 inst_cellmath__48_I29657 (.Y(N23273), .A(N7812));
INVX2 inst_cellmath__48_I29658 (.Y(N23275), .A(N23273));
CLKXOR2X1 inst_cellmath__48_I29659 (.Y(N45499), .A(N45494), .B(N23275));
CLKINVX4 inst_cellmath__48_I29660 (.Y(N10973), .A(N45499));
INVXL buf1_A_I30577 (.Y(N45771), .A(N45499));
INVXL buf1_A_I30578 (.Y(inst_cellmath__61[11]), .A(N45771));
NAND2XL inst_cellmath__48_I29449 (.Y(N44986), .A(N7395), .B(N7525));
NOR2XL inst_cellmath__48_I29450 (.Y(N707), .A(N44986), .B(inst_cellmath__42[5]));
MXI2XL inst_cellmath__48_I1361 (.Y(N7390), .A(N7335), .B(N7464), .S0(N7395));
MXI2XL inst_cellmath__48_I1362 (.Y(N7446), .A(N7392), .B(N7518), .S0(N7395));
MXI2XL inst_cellmath__48_I1363 (.Y(N7498), .A(N7448), .B(N7320), .S0(N7395));
MXI2XL inst_cellmath__48_I1364 (.Y(N7555), .A(N7501), .B(N7375), .S0(N7395));
MXI2XL inst_cellmath__48_I1365 (.Y(N7355), .A(N7557), .B(N7434), .S0(N7395));
MXI2X1 inst_cellmath__48_I1366 (.Y(N7412), .A(N7357), .B(N7487), .S0(N7395));
MXI2X1 inst_cellmath__48_I1367 (.Y(N7469), .A(N7414), .B(N7544), .S0(N7395));
MXI2X1 inst_cellmath__48_I1368 (.Y(N7524), .A(N7525), .B(N7343), .S0(N7395));
MXI2XL inst_cellmath__48_I1369 (.Y(N7324), .A(N7381), .B(N7400), .S0(N7395));
MXI2X1 inst_cellmath__48_I1370 (.Y(N7379), .A(N7492), .B(N7456), .S0(N7395));
MXI2XL inst_cellmath__48_I1371 (.Y(N7438), .A(N7349), .B(N7510), .S0(N7395));
MXI2XL inst_cellmath__48_I1373 (.Y(N7549), .A(N7570), .B(N7366), .S0(N7395));
MXI2XL inst_cellmath__48_I1374 (.Y(N7348), .A(N7428), .B(N7423), .S0(N7395));
NAND2XL inst_cellmath__48_I1375 (.Y(N7404), .A(N7395), .B(N7477));
NAND2XL inst_cellmath__48_I1376 (.Y(N7513), .A(N7395), .B(N7535));
NAND2XL inst_cellmath__48_I1377 (.Y(N7370), .A(N7395), .B(N7335));
NAND2XL inst_cellmath__48_I1378 (.Y(N7480), .A(N7395), .B(N7392));
NAND2XL inst_cellmath__48_I1379 (.Y(N7337), .A(N7395), .B(N7448));
NAND2X1 inst_cellmath__48_I1380 (.Y(N7450), .A(N7395), .B(N7501));
NAND2XL inst_cellmath__48_I1381 (.Y(N7559), .A(N7395), .B(N7557));
NAND2XL inst_cellmath__48_I1382 (.Y(N7416), .A(N7395), .B(N7357));
NAND2XL inst_cellmath__48_I1383 (.Y(N7528), .A(N7414), .B(N7395));
NAND2XL inst_cellmath__48_I1385 (.Y(N7494), .A(N7395), .B(N7381));
NOR2XL inst_cellmath__48_I1394 (.Y(N684), .A(inst_cellmath__42[5]), .B(N7390));
NOR2XL inst_cellmath__48_I1395 (.Y(N685), .A(inst_cellmath__42[5]), .B(N7446));
NOR2X1 inst_cellmath__48_I1396 (.Y(N686), .A(inst_cellmath__42[5]), .B(N7498));
NOR2XL inst_cellmath__48_I1397 (.Y(N687), .A(inst_cellmath__42[5]), .B(N7555));
NOR2XL inst_cellmath__48_I1398 (.Y(N688), .A(inst_cellmath__42[5]), .B(N7355));
NOR2X1 inst_cellmath__48_I1399 (.Y(N689), .A(inst_cellmath__42[5]), .B(N7412));
NOR2X1 inst_cellmath__48_I1400 (.Y(N690), .A(inst_cellmath__42[5]), .B(N7469));
NOR2X2 inst_cellmath__48_I1401 (.Y(N691), .A(inst_cellmath__42[5]), .B(N7524));
NOR2XL inst_cellmath__48_I1402 (.Y(N692), .A(inst_cellmath__42[5]), .B(N7324));
NOR2X2 inst_cellmath__48_I1403 (.Y(N693), .A(inst_cellmath__42[5]), .B(N7379));
NOR2XL inst_cellmath__48_I1404 (.Y(N694), .A(inst_cellmath__42[5]), .B(N7438));
NOR2XL inst_cellmath__48_I1406 (.Y(N696), .A(inst_cellmath__42[5]), .B(N7549));
NOR2XL inst_cellmath__48_I1407 (.Y(N697), .A(inst_cellmath__42[5]), .B(N7348));
NOR2X1 inst_cellmath__48_I1408 (.Y(N698), .A(inst_cellmath__42[5]), .B(N7404));
NOR2X1 inst_cellmath__48_I1409 (.Y(N699), .A(inst_cellmath__42[5]), .B(N7513));
NOR2XL inst_cellmath__48_I1410 (.Y(N700), .A(inst_cellmath__42[5]), .B(N7370));
NOR2XL inst_cellmath__48_I1411 (.Y(N701), .A(inst_cellmath__42[5]), .B(N7480));
NOR2X1 inst_cellmath__48_I1412 (.Y(N702), .A(inst_cellmath__42[5]), .B(N7337));
NOR2X1 inst_cellmath__48_I1413 (.Y(N703), .A(inst_cellmath__42[5]), .B(N7450));
NOR2XL inst_cellmath__48_I1414 (.Y(N704), .A(inst_cellmath__42[5]), .B(N7559));
NOR2XL inst_cellmath__48_I1415 (.Y(N705), .A(inst_cellmath__42[5]), .B(N7416));
NOR2XL inst_cellmath__48_I1416 (.Y(N706), .A(inst_cellmath__42[5]), .B(N7528));
NOR2XL inst_cellmath__48_I1418 (.Y(N708), .A(N7494), .B(inst_cellmath__42[5]));
XOR2XL cynw_cm_float_cos_I1420 (.Y(N493), .A(N708), .B(N707));
INVX1 inst_cellmath__61_0_I1422 (.Y(N7809), .A(N691));
INVX1 inst_cellmath__61_0_I1423 (.Y(N7833), .A(N693));
INVXL inst_cellmath__61_0_I10573 (.Y(N23278), .A(N23273));
INVX2 inst_cellmath__61_0_I10572 (.Y(N23277), .A(N23273));
INVX2 inst_cellmath__61_0_I10571 (.Y(N23276), .A(N23273));
INVX2 inst_cellmath__61_0_I10569 (.Y(N23274), .A(N23273));
CLKXOR2X1 inst_cellmath__61_0_I11191 (.Y(inst_cellmath__61[0]), .A(N684), .B(N23278));
CLKXOR2X1 inst_cellmath__61_0_I1430 (.Y(inst_cellmath__61[1]), .A(N685), .B(N23278));
XOR2X4 inst_cellmath__61_0_I10831 (.Y(inst_cellmath__61[2]), .A(N23277), .B(N686));
CLKXOR2X1 inst_cellmath__61_0_I1432 (.Y(inst_cellmath__61[3]), .A(N23274), .B(N687));
CLKXOR2X1 inst_cellmath__61_0_I1433 (.Y(inst_cellmath__61[4]), .A(N23274), .B(N688));
CLKXOR2X1 inst_cellmath__61_0_I1434 (.Y(inst_cellmath__61[5]), .A(N689), .B(N23274));
XNOR2X1 inst_cellmath__61_0_I1435 (.Y(inst_cellmath__61[6]), .A(N7812), .B(N690));
MXI2X1 inst_cellmath__61_0_I1436 (.Y(inst_cellmath__61[7]), .A(N7809), .B(N691), .S0(N23274));
XOR2X1 inst_cellmath__61_0_I1437 (.Y(inst_cellmath__61[8]), .A(N692), .B(N23274));
MXI2X1 inst_cellmath__61_0_I1438 (.Y(inst_cellmath__61[9]), .A(N7833), .B(N693), .S0(N23275));
CLKXOR2X1 inst_cellmath__61_0_I1439 (.Y(inst_cellmath__61[10]), .A(N694), .B(N23275));
CLKXOR2X1 inst_cellmath__61_0_I1441 (.Y(inst_cellmath__61[12]), .A(N696), .B(N23275));
XOR2X1 inst_cellmath__61_0_I1442 (.Y(inst_cellmath__61[13]), .A(N697), .B(N23276));
CLKXOR2X1 inst_cellmath__61_0_I1443 (.Y(inst_cellmath__61[14]), .A(N23277), .B(N698));
CLKXOR2X1 inst_cellmath__61_0_I1444 (.Y(inst_cellmath__61[15]), .A(N699), .B(N23277));
CLKXOR2X1 inst_cellmath__61_0_I1445 (.Y(inst_cellmath__61[16]), .A(N700), .B(N23277));
CLKXOR2X1 inst_cellmath__61_0_I1446 (.Y(inst_cellmath__61[17]), .A(N701), .B(N23277));
CLKXOR2X1 inst_cellmath__61_0_I1447 (.Y(inst_cellmath__61[18]), .A(N702), .B(N23275));
CLKXOR2X1 inst_cellmath__61_0_I1448 (.Y(inst_cellmath__61[19]), .A(N703), .B(N23276));
CLKXOR2X1 inst_cellmath__61_0_I1449 (.Y(inst_cellmath__61[20]), .A(N704), .B(N23276));
CLKXOR2X1 inst_cellmath__61_0_I1450 (.Y(inst_cellmath__61[21]), .A(N705), .B(N23276));
CLKXOR2X1 inst_cellmath__61_0_I1451 (.Y(inst_cellmath__61[22]), .A(N706), .B(N23276));
INVX3 cynw_cm_float_cos_I361 (.Y(N3808), .A(inst_cellmath__61[6]));
CLKINVX4 cynw_cm_float_cos_I362 (.Y(N3809), .A(inst_cellmath__61[10]));
INVX1 cynw_cm_float_cos_I363 (.Y(N3810), .A(N3809));
INVX2 cynw_cm_float_cos_I5 (.Y(inst_cellmath__115__W1[0]), .A(inst_cellmath__61[16]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1454 (.Y(N8330), .A(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1455 (.Y(N8985), .A(inst_cellmath__61[20]), .B(inst_cellmath__61[21]));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I11197 (.Y(N7912), .A(N8330), .B(N8985));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1459 (.Y(N8703), .A(inst_cellmath__61[19]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1460 (.Y(N8536), .A(inst_cellmath__61[17]), .B(inst_cellmath__61[18]));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10838 (.Y(N8289), .A(N8703), .B(N8536));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1464 (.Y(N8463), .A(N8289), .B(N7912));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1465 (.Y(N8122), .A(inst_cellmath__61[17]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1466 (.Y(N8375), .A(inst_cellmath__61[18]), .B(N8122));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1467 (.Y(N9127), .A(N8375), .B(N8703));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1468 (.Y(N8396), .A(N9127));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1470 (.Y(N8309), .A(N7912), .B(N8396));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1471 (.Y(N7949), .A(inst_cellmath__61[18]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1472 (.Y(N8231), .A(inst_cellmath__61[17]), .B(N7949));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10840 (.Y(N8511), .A(N8703), .B(N8231));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1476 (.Y(N8756), .A(N7912), .B(N8511));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1477 (.Y(N9050), .A(N8122), .B(N7949));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1478 (.Y(N8780), .A(N9050), .B(N8703));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1479 (.Y(N8083), .A(N8780));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1481 (.Y(N8333), .A(N7912), .B(N8083));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10692 (.Y(N8206), .A(inst_cellmath__61[19]), .B(N8536));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1485 (.Y(N7999), .A(N7912), .B(N8206));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1486 (.Y(N9026), .A(N8375), .B(inst_cellmath__61[19]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1487 (.Y(N8306), .A(N9026));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1489 (.Y(N8185), .A(N7912), .B(N8306));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I11201 (.Y(N7888), .A(inst_cellmath__61[19]), .B(N8231));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1493 (.Y(N8705), .A(N7912), .B(N7888));
AND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1494 (.Y(N8161), .A(N9050), .B(inst_cellmath__61[19]));
INVX2 inst_cellmath__195__80__2WWMM_2WWMM_I1495 (.Y(N8676), .A(N8161));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1497 (.Y(N8928), .A(N7912), .B(N8676));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1498 (.Y(N8291), .A(inst_cellmath__61[20]));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1499 (.Y(N8554), .A(inst_cellmath__61[21]), .B(N8291));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I11306 (.Y(N8804), .A(N8330), .B(N8554));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1503 (.Y(N9132), .A(N8289), .B(N8804));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1504 (.Y(N8146), .A(N8804), .B(N8396));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1505 (.Y(N8399), .A(N8804), .B(N8511));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1506 (.Y(N8654), .A(N8804), .B(N8083));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1507 (.Y(N8949), .A(N8804), .B(N8206));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1508 (.Y(N7976), .A(N8804), .B(N8306));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1509 (.Y(N8753), .A(N8804), .B(N7888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1510 (.Y(N8513), .A(N8804), .B(N8676));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1511 (.Y(N8782), .A(inst_cellmath__61[21]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1512 (.Y(N9075), .A(inst_cellmath__61[20]), .B(N8782));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10846 (.Y(N8923), .A(N8330), .B(N9075));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1516 (.Y(N8351), .A(N8289), .B(N8923));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1517 (.Y(N8615), .A(N8923), .B(N8396));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1518 (.Y(N8904), .A(N8511), .B(N8923));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1519 (.Y(N8598), .A(N8923), .B(N8083));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1520 (.Y(N7911), .A(N8923), .B(N8206));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1521 (.Y(N8462), .A(N8923), .B(N8306));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1522 (.Y(N8441), .A(N8923), .B(N7888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1523 (.Y(N9028), .A(N8923), .B(N8676));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1524 (.Y(N8037), .A(N8291), .B(N8782));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I11204 (.Y(N7905), .A(N8330), .B(N8037));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1528 (.Y(N8575), .A(N8289), .B(N7905));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1529 (.Y(N8853), .A(N8396), .B(N7905));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1530 (.Y(N8288), .A(N8511), .B(N7905));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1531 (.Y(N8164), .A(N7905), .B(N8083));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1532 (.Y(N8419), .A(N7905), .B(N8206));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1533 (.Y(N8677), .A(N7905), .B(N8306));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1534 (.Y(N8977), .A(N7905), .B(N7888));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1535 (.Y(N7995), .A(N7905), .B(N8676));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10848 (.Y(N8010), .A(inst_cellmath__61[22]), .B(N8985));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1539 (.Y(N8532), .A(N8289), .B(N8010));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1540 (.Y(N8806), .A(N8010), .B(N8396));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1541 (.Y(N9101), .A(N8010), .B(N8511));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1542 (.Y(N8112), .A(N8010), .B(N8083));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1543 (.Y(N8370), .A(N8010), .B(N8206));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1544 (.Y(N8633), .A(N8010), .B(N8306));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1545 (.Y(N8925), .A(N8010), .B(N7888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1546 (.Y(N7943), .A(N8010), .B(N8676));
NAND2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10849 (.Y(N8828), .A(N8554), .B(inst_cellmath__61[22]));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1550 (.Y(N8483), .A(N8289), .B(N8828));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1551 (.Y(N8748), .A(N8828), .B(N8396));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1552 (.Y(N9046), .A(N8828), .B(N8511));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1553 (.Y(N8057), .A(N8828), .B(N8083));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1554 (.Y(N8323), .A(N8828), .B(N8206));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1555 (.Y(N8595), .A(N8828), .B(N8306));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1556 (.Y(N8875), .A(N8828), .B(N7888));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1557 (.Y(N7907), .A(N8828), .B(N8676));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I11205 (.Y(N8389), .A(inst_cellmath__61[22]), .B(N9075));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1561 (.Y(N7971), .A(N8289), .B(N8389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1562 (.Y(N8701), .A(N8396), .B(N8389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1563 (.Y(N9003), .A(N8389), .B(N8511));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1564 (.Y(N8011), .A(N8083), .B(N8389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1565 (.Y(N8286), .A(N8206), .B(N8389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1566 (.Y(N8548), .A(N8306), .B(N8389));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1567 (.Y(N8831), .A(N8389), .B(N7888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1568 (.Y(N9123), .A(N8389), .B(N8676));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I11307 (.Y(N8506), .A(inst_cellmath__61[22]), .B(N8037));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1572 (.Y(N8392), .A(N8289), .B(N8506));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1573 (.Y(N8651), .A(N8396), .B(N8506));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1574 (.Y(N9071), .A(N8511), .B(N8506));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1575 (.Y(N7967), .A(N8506), .B(N8083));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I10703 (.Y(N8609), .A(N8206), .B(N8506));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1579 (.Y(N8901), .A(N8506), .B(N8306));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1580 (.Y(N8773), .A(N8506), .B(N7888));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1581 (.Y(N9066), .A(N8506), .B(N8676));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1582 (.Y(N8201), .A(N8463));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1583 (.Y(N8457), .A(N8309));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1584 (.Y(N8205), .A(N8309), .B(N8463));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1585 (.Y(N8569), .A(N8756));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1586 (.Y(N8847), .A(N8333));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1587 (.Y(N8724), .A(N8756), .B(N8333));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1588 (.Y(N8035), .A(N7999), .B(N8185));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1589 (.Y(N8799), .A(N8185));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1590 (.Y(N9092), .A(N7999));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1591 (.Y(N8104), .A(N8705));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1592 (.Y(N8363), .A(N8928));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1593 (.Y(N8572), .A(N8705), .B(N8928));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1594 (.Y(N7887), .A(N8146), .B(N9132));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1595 (.Y(N8049), .A(N9132));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1596 (.Y(N8587), .A(N8146));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1597 (.Y(N8416), .A(N8399), .B(N8654));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1598 (.Y(N8434), .A(N8654));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1599 (.Y(N8692), .A(N8399));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1600 (.Y(N8997), .A(N7976));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1601 (.Y(N8825), .A(N8949));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I11308 (.Y(N8646), .A(N7976), .B(N8949));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1607 (.Y(N8762), .A(N8753));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I11208 (.Y(N8603), .A(N8753), .B(N8513));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1612 (.Y(N8890), .A(N8513));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1613 (.Y(N7919), .A(N8351));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1614 (.Y(N8195), .A(N8351), .B(N8615));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1615 (.Y(N8713), .A(N8195));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1617 (.Y(N9140), .A(N8615));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1618 (.Y(N8154), .A(N8598));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1619 (.Y(N8109), .A(N8598), .B(N8904));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1620 (.Y(N8962), .A(N8904));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1621 (.Y(N8628), .A(N8462), .B(N7911));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1622 (.Y(N8520), .A(N7911));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1623 (.Y(N8795), .A(N8462));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1624 (.Y(N9086), .A(N9028));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1625 (.Y(N8097), .A(N8441));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1626 (.Y(N8912), .A(N8441), .B(N9028));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1627 (.Y(N9034), .A(N8853));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1629 (.Y(N8043), .A(N8575));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1630 (.Y(N8481), .A(N8853), .B(N8575));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1631 (.Y(N8859), .A(N8164));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1632 (.Y(N9044), .A(N8288), .B(N8164));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1633 (.Y(N8427), .A(N8288));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1634 (.Y(N8320), .A(N8677), .B(N8419));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1635 (.Y(N8001), .A(N8677));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1636 (.Y(N8274), .A(N8419));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1637 (.Y(N8870), .A(N7995), .B(N8977));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1638 (.Y(N9109), .A(N8977));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1639 (.Y(N8125), .A(N7995));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1640 (.Y(N8178), .A(N8532), .B(N8806));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1641 (.Y(N8931), .A(N8532));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1642 (.Y(N9052), .A(N8806));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1644 (.Y(N8066), .A(N8112));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1645 (.Y(N8187), .A(N9101));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1646 (.Y(N8697), .A(N9101), .B(N8112));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1647 (.Y(N9012), .A(N8370));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I10706 (.Y(N8837), .A(N8633), .B(N8370));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1651 (.Y(N9134), .A(N8633));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1652 (.Y(N8545), .A(N7943), .B(N8925));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1653 (.Y(N8659), .A(N7943));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1654 (.Y(N8953), .A(N8925));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1655 (.Y(N7978), .A(N8483));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1656 (.Y(N9119), .A(N8483), .B(N8748));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1657 (.Y(N8785), .A(N8748));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1658 (.Y(N9077), .A(N8057));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1659 (.Y(N8207), .A(N9046));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1661 (.Y(N8725), .A(N8057), .B(N9046));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1662 (.Y(N9029), .A(N8323));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1663 (.Y(N8039), .A(N8595));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1664 (.Y(N8943), .A(N8595), .B(N8323));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1665 (.Y(N8854), .A(N7907));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1666 (.Y(N8166), .A(N7907), .B(N8875));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1667 (.Y(N8421), .A(N8875));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1668 (.Y(N8680), .A(N8701));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1669 (.Y(N8770), .A(N7971), .B(N8701));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1670 (.Y(N8269), .A(N7971));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1671 (.Y(N8077), .A(N8011), .B(N9003));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1672 (.Y(N9103), .A(N8011));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1673 (.Y(N8116), .A(N9003));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1674 (.Y(N8608), .A(N8548), .B(N8286));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1675 (.Y(N8927), .A(N8286));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1676 (.Y(N7945), .A(N8548));
OR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1677 (.Y(N8227), .A(N8831), .B(N9123));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1678 (.Y(N8750), .A(N8227));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1680 (.Y(N8876), .A(N9123));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1681 (.Y(N7908), .A(N8831));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1682 (.Y(N8181), .A(N8392));
NOR2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1683 (.Y(N8456), .A(N8392), .B(N8651));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1684 (.Y(N9004), .A(N8651));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1685 (.Y(N9022), .A(N9071), .B(N7967));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1686 (.Y(N8550), .A(N9071));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1687 (.Y(N8832), .A(N7967));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1688 (.Y(N9125), .A(N8901));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I1689 (.Y(N8304), .A(N8901), .B(N8609));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1690 (.Y(N8653), .A(N8609));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1691 (.Y(N8947), .A(N9066));
NOR2X2 inst_cellmath__195__80__2WWMM_2WWMM_I10707 (.Y(N8776), .A(N9066), .B(N8773));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1695 (.Y(N9069), .A(N8773));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1696 (.Y(N8216), .A(N9012), .B(N7919));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1697 (.Y(N8006), .A(N7978), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1698 (.Y(N8280), .A(N9034), .B(N8628));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1699 (.Y(N8159), .A(N8035), .B(N8178));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1700 (.Y(N8826), .A(N8066), .B(N9077));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1701 (.Y(N9117), .A(N9086), .B(N8569));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1702 (.Y(N8136), .A(N7887), .B(N8762));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1703 (.Y(N7921), .A(N8201), .B(N8859));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1704 (.Y(N8130), .A(N8416), .B(N8750));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1705 (.Y(N8606), .A(N8870), .B(N9022));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1706 (.Y(N8715), .A(N8077), .B(N8216));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1707 (.Y(N8766), .A(N9125), .B(N9029), .C(N8006));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1708 (.Y(N9060), .A(N8280), .B(N8826));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1709 (.Y(N8073), .A(N9117), .B(N8159));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1710 (.Y(N8344), .A(N8136), .B(N8130));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1711 (.Y(N8197), .A(N7921), .B(N9060));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1712 (.Y(N8452), .A(N8073), .B(N8344));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1713 (.Y(N9019), .A(N8715), .B(N8452));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1714 (.Y(N8033), .A(N8606), .B(N8766), .C(N8197));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1716 (.Y(N8666), .A(N8931), .B(N7919));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1717 (.Y(N8964), .A(N8043), .B(N8181));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1718 (.Y(N7986), .A(N8520), .B(N9125));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1719 (.Y(N8613), .A(N8320), .B(N8608));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1720 (.Y(N8899), .A(N8613));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1721 (.Y(N7990), .A(N9086), .B(N8770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1722 (.Y(N8099), .A(N8847), .B(N9119));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1723 (.Y(N7923), .A(N8154), .B(N8859));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1724 (.Y(N8622), .A(N8603));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1725 (.Y(N8914), .A(N8622), .B(N8964));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1726 (.Y(N8721), .A(N8545));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1727 (.Y(N8199), .A(N8049), .B(N8039));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1728 (.Y(N8469), .A(N8721), .B(N8199));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1729 (.Y(N8735), .A(N8666), .B(N7986));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1730 (.Y(N9037), .A(N8099), .B(N8899));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1731 (.Y(N8312), .A(N7923), .B(N8606));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1732 (.Y(N8862), .A(N8914), .B(N8469));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1733 (.Y(N8420), .A(N9077), .B(N8312), .C(N8104));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1734 (.Y(N8429), .A(N7990), .B(N8420));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1735 (.Y(N8845), .A(N8735), .B(N9037));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1736 (.Y(N8172), .A(N8862), .B(N8845));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1738 (.Y(N8523), .A(N8320), .B(N8628));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1739 (.Y(N9091), .AN(N8195), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1740 (.Y(N8934), .A(N8066), .B(N8434));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1741 (.Y(N8362), .A(N8943), .B(N8837));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1742 (.Y(N8233), .A(N8876), .B(N8847));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1743 (.Y(N8491), .A(N7887), .B(N8481));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1744 (.Y(N8758), .A(N9119), .B(N9109));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1745 (.Y(N8643), .A(N8207), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1747 (.Y(N8336), .A(N8109), .B(N9044));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1748 (.Y(N8884), .A(N9091), .B(N8362));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1749 (.Y(N7915), .A(N8233), .B(N8934));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1750 (.Y(N8191), .A(N8523), .B(N8491));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1751 (.Y(N8445), .A(N8758), .B(N8336));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29767 (.Y(N9015), .A(N8659), .B(N9022), .C(N8304), .D(N8643));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1754 (.Y(N8295), .A(N8191), .B(N8445));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1755 (.Y(N8916), .A(N8884), .B(N7915));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1756 (.Y(N8560), .A(N8295), .B(N8916));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1758 (.Y(N8251), .A(N9125), .B(N8001));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1759 (.Y(N8517), .A(N8795), .B(N9140));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1760 (.Y(N8788), .A(N8799), .B(N9052));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1761 (.Y(N9080), .A(N8039), .B(N9134));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1762 (.Y(N8090), .A(N8680), .B(N9034));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1763 (.Y(N8355), .A(N8608), .B(N9077));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1764 (.Y(N8917), .A(N9086), .B(N8876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1765 (.Y(N8908), .A(N8187), .B(N8947));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1766 (.Y(N7933), .A(N8854), .B(N8659));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1767 (.Y(N8209), .A(N8762), .B(N8416));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1768 (.Y(N8464), .A(N8517), .B(N8788));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1769 (.Y(N8672), .A(N9044));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1770 (.Y(N8423), .A(N8917), .B(N9080));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1771 (.Y(N8272), .A(N8423), .B(N8464));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1772 (.Y(N8682), .A(N8090), .B(N8908));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1773 (.Y(N8856), .A(N8251), .B(N7933));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1774 (.Y(N7892), .A(N8355), .B(N8209));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1775 (.Y(N8983), .A(N8181), .B(N9022), .C(N8682));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1776 (.Y(N8811), .A(N8856), .B(N7892));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1777 (.Y(N8120), .A(N8272), .B(N8672));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1778 (.Y(N9106), .A(N8811), .B(N8983));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1780 (.Y(N8182), .A(N8997), .B(N8795));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1781 (.Y(N8398), .A(N8481), .B(N7908));
INVX1 inst_cellmath__195__80__2WWMM_2WWMM_I1782 (.Y(N8970), .A(N8572));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1783 (.Y(N8315), .A(N8274), .B(N8049));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1784 (.Y(N9128), .A(N8970), .B(N8315));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1785 (.Y(N8781), .A(N8288), .B(N7999), .C(N8398));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1786 (.Y(N8247), .A(N9077), .B(N8550), .C(N8870), .D(N8943));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1787 (.Y(N7973), .A(N8182), .B(N8006), .C(N9128));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1788 (.Y(N8512), .A(N8247), .B(N7973));
NAND2BXL inst_cellmath__195__80__2WWMM_2WWMM_I1790 (.Y(N8219), .AN(N9132), .B(N8825));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1791 (.Y(N8142), .A(N8927), .B(N9004));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1792 (.Y(N8741), .A(N8799), .B(N8039));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1793 (.Y(N8574), .A(N8713), .B(N8066));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1794 (.Y(N8851), .A(N7908), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1795 (.Y(N7948), .A(N9103), .B(N8550));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1796 (.Y(N8162), .A(N8762), .B(N8776));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1797 (.Y(N8530), .A(N8545), .B(N8109));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1798 (.Y(N8973), .A(N8741), .B(N7948));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1799 (.Y(N7994), .A(N8851), .B(N8574));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1800 (.Y(N8110), .AN(N8162), .B(N8320), .C(N9034));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1801 (.Y(N8630), .A(N8142), .B(N8219), .C(N8530));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1802 (.Y(N9099), .A(N8973), .B(N7994));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1803 (.Y(N8368), .A(N8110), .B(N9099));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1805 (.Y(N8056), .A(N9092), .B(N8181));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1806 (.Y(N8321), .A(N8274), .B(N8795));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1807 (.Y(N8592), .A(N8927), .B(N9052));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1808 (.Y(N8873), .A(N8039), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1809 (.Y(N9020), .A(N8785), .B(N8646));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1810 (.Y(N8179), .A(N8713), .B(N8692));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1811 (.Y(N8439), .A(N8953), .B(N8847));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1812 (.Y(N8685), .A(N8854), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1813 (.Y(N8048), .A(N8125), .B(N8832));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1814 (.Y(N8829), .A(N8603), .B(N8572));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1815 (.Y(N8365), .A(N8109));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1816 (.Y(N8507), .A(N8592), .B(N8056));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1817 (.Y(N8648), .A(N8048), .B(N8321));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1818 (.Y(N8944), .A(N8908), .B(N8439));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1819 (.Y(N7965), .A(N8685), .B(N8873));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1820 (.Y(N8241), .A(N8179), .B(N8829));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1821 (.Y(N8771), .A(N8507), .B(N7921));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1822 (.Y(N9063), .A(N8648), .B(N8944));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1823 (.Y(N8896), .A(N7965), .B(N8241));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1824 (.Y(N8202), .A(N9020), .B(N8365), .C(N9063));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1825 (.Y(N7924), .A(N8896), .B(N8771));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1827 (.Y(N8967), .A(N8713), .B(N8178));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1828 (.Y(N7991), .A(N9077), .B(N8837));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1829 (.Y(N8261), .A(N8569), .B(N7887));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1830 (.Y(N8525), .A(N8481), .B(N8890));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1831 (.Y(N8801), .A(N8550), .B(N8697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1832 (.Y(N9093), .A(N8416), .B(N8776));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1833 (.Y(N8220), .A(N8261), .B(N8801));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1834 (.Y(N8474), .A(N8741), .B(N8525));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1835 (.Y(N7902), .A(N8427), .B(N8646), .C(N8220), .D(N8474));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I1838 (.Y(N8435), .AN(N8463), .B(N8545), .C(N8166), .D(N8870));
OR4XL inst_cellmath__195__80__2WWMM_2WWMM_I29800 (.Y(N8865), .A(N7991), .B(N9093), .C(N8967), .D(N8899));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1840 (.Y(N8175), .A(N7902), .B(N8365));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1841 (.Y(N8694), .A(N8435), .B(N8865));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1843 (.Y(N8626), .A(N8457), .B(N9092));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1844 (.Y(N8135), .A(N8997), .B(N7978));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1845 (.Y(N8386), .A(N9052), .B(N8039));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1846 (.Y(N8647), .A(N9134), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1847 (.Y(N8939), .A(N8587), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1848 (.Y(N8236), .A(N8628), .B(N8569));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1849 (.Y(N8497), .A(N8187), .B(N8854));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1850 (.Y(N8764), .A(N8207), .B(N8550));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1851 (.Y(N7940), .A(N8750), .B(N8776));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1852 (.Y(N8342), .A(N8622), .B(N8939));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1853 (.Y(N8891), .A(N8626), .B(N8870));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1854 (.Y(N8196), .A(N8721), .B(N8135));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1855 (.Y(N9017), .A(N8497), .B(N8236));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1856 (.Y(N8030), .A(N8647), .B(N8764));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1857 (.Y(N8300), .A(N7940), .B(N8386));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1858 (.Y(N8564), .A(N8899), .B(N8891));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1859 (.Y(N8842), .A(N9017), .B(N8030));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1860 (.Y(N9141), .A(N8342), .B(N8300));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1861 (.Y(N8155), .A(N8196), .B(N8564));
NOR4BBX1 inst_cellmath__195__80__2WWMM_2WWMM_I1862 (.Y(N8665), .AN(N8181), .BN(N9125), .C(N8365), .D(N8842));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1863 (.Y(N8963), .A(N9141), .B(N8155));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1865 (.Y(N8796), .A(N8931), .B(N8043));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1866 (.Y(N8096), .A(N8785), .B(N8587));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1867 (.Y(N8620), .A(N8205), .B(N8646));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1868 (.Y(N8276), .A(N8608), .B(N8713));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1869 (.Y(N8214), .A(N8421), .B(N8770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1870 (.Y(N8467), .A(N8569), .B(N8187));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1871 (.Y(N8732), .A(N9109), .B(N8890));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1872 (.Y(N8044), .A(N8659), .B(N8859));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1873 (.Y(N8433), .A(N8416), .B(N8912));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1874 (.Y(N8987), .A(N8796), .B(N8096));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1875 (.Y(N8816), .A(N9022), .B(N8077));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1876 (.Y(N7897), .A(N8214), .B(N8732));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1877 (.Y(N8994), .A(N8799), .B(N9134));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1878 (.Y(N8170), .A(N8620), .B(N8994));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1879 (.Y(N8428), .A(N8001), .B(N8962), .C(N8943), .D(N8181));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1880 (.Y(N8686), .A(N8467), .B(N8044));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1881 (.Y(N8275), .A(N8276), .B(N8433));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1882 (.Y(N8126), .A(N8686), .B(N8275));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I1883 (.Y(N7951), .A(N7897), .B(N8987), .C(N8643), .D(N8170));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1884 (.Y(N8932), .A(N8428), .B(N8816), .C(N8126));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1886 (.Y(N8995), .A(N9052), .B(N9134));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1887 (.Y(N8188), .A(N9034), .B(N8785));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1888 (.Y(N8706), .A(N8035), .B(N8066));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1889 (.Y(N9013), .A(N8434), .B(N8847));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1890 (.Y(N8021), .A(N7887), .B(N7908));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1891 (.Y(N8293), .A(N8947), .B(N8659));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1892 (.Y(N8279), .A(N9103), .B(N8762));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1893 (.Y(N9135), .A(N8725), .B(N8166));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1894 (.Y(N8515), .A(N9004), .B(N9029), .C(N8182));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1895 (.Y(N8402), .A(N8995), .B(N8901));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1896 (.Y(N8660), .A(N8188), .B(N9135));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1899 (.Y(N9079), .A(N8402), .B(N8660));
OR4XL inst_cellmath__195__80__2WWMM_2WWMM_I29816 (.Y(N8906), .A(N8706), .B(N9013), .C(N8293), .D(N8279));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1901 (.Y(N8208), .A(N8021), .B(N7923), .C(N9079));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1902 (.Y(N7932), .A(N8515), .B(N8899), .C(N8906));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1904 (.Y(N8751), .A(N9034), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1905 (.Y(N8981), .A(N8608), .B(N8628));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1906 (.Y(N7997), .A(N8692), .B(N8837));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1907 (.Y(N8270), .A(N8569), .B(N9119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1908 (.Y(N8809), .A(N8363), .B(N8659));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1909 (.Y(N9104), .A(N8859), .B(N8697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1910 (.Y(N8117), .A(N8725), .B(N8750));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1911 (.Y(N8824), .A(N8166), .B(N8776));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1912 (.Y(N7946), .A(N8931), .B(N8457), .C(N8109));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1913 (.Y(N9005), .A(N7971), .B(N8751), .C(N8651));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1914 (.Y(N8060), .A(N8809), .B(N8270));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1915 (.Y(N8327), .A(N8741), .B(N8824));
NAND4BBXL inst_cellmath__195__80__2WWMM_2WWMM_I1916 (.Y(N8877), .AN(N8219), .BN(N8048), .C(N8603), .D(N8077));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1917 (.Y(N7909), .A(N9104));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1918 (.Y(N8551), .AN(N7909), .B(N7997), .C(N8117));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1919 (.Y(N8440), .A(N8981), .B(N7946));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1920 (.Y(N8014), .A(N9005), .B(N8440));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1921 (.Y(N8382), .A(N8060), .B(N8327));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1922 (.Y(N8287), .A(N8877), .B(N8382));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1923 (.Y(N753), .AN(N8014), .B(N8551), .C(N8287));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1924 (.Y(N8777), .A(N8274), .B(N8927));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1925 (.Y(N9070), .A(N8785), .B(N8304));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1926 (.Y(N8132), .A(N8178), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1927 (.Y(N8055), .A(N8847), .B(N8481));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1928 (.Y(N8203), .A(N7908), .B(N8762));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1929 (.Y(N8722), .A(N8598), .B(N8777));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1930 (.Y(N8264), .A(N8870), .B(N8626));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1931 (.Y(N9055), .A(N8692), .B(N8953));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1932 (.Y(N8673), .A(N9055), .B(N8132));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1933 (.Y(N8849), .A(N9070), .B(N8203));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1934 (.Y(N7885), .A(N8055), .B(N8826));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1935 (.Y(N8415), .A(N8116), .B(N8713), .C(N8722));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1936 (.Y(N8972), .A(N8859), .B(N8776), .C(N8673));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1937 (.Y(N8803), .A(N8849), .B(N7885));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1938 (.Y(N8108), .A(N8264), .B(N8415));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1939 (.Y(N9096), .A(N8803), .B(N8972));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1941 (.Y(N8645), .A(N8825), .B(N8795));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1942 (.Y(N8868), .A(N8269), .B(N8320));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1943 (.Y(N8544), .A(N8962), .B(N8421));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1944 (.Y(N8281), .A(N8125), .B(N9103));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1945 (.Y(N8076), .A(N8592), .B(N8917));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1946 (.Y(N8534), .A(N8572), .B(N8545));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I1947 (.Y(N7963), .A(N9029), .B(N7978), .C(N8626));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1948 (.Y(N8941), .A(N8525), .B(N8261));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1949 (.Y(N8238), .A(N7963), .B(N8534));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1950 (.Y(N8504), .A(N8868), .B(N7991));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I1951 (.Y(N9061), .A(N8281), .B(N8645), .C(N9091));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1952 (.Y(N7922), .AN(N8544), .B(N8076), .C(N8859));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1953 (.Y(N8607), .A(N8941), .B(N8504));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1954 (.Y(N8200), .A(N7922), .B(N8607));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1956 (.Y(N8846), .A(N8201), .B(N8653));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1957 (.Y(N7882), .A(N8043), .B(N8274));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1958 (.Y(N8668), .A(N8116), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1959 (.Y(N8966), .A(N8608), .B(N8035));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1960 (.Y(N7989), .A(N8434), .B(N9069));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1961 (.Y(N8259), .A(N8837), .B(N8876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1962 (.Y(N8522), .A(N9119), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1963 (.Y(N8798), .A(N8363), .B(N8550));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1964 (.Y(N9089), .A(N8697), .B(N8166));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1965 (.Y(N8101), .A(N8846), .B(N7882));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I1966 (.Y(N7937), .AN(N8721), .B(N8587), .C(N9004));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1967 (.Y(N8218), .A(N7989), .B(N8645));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1968 (.Y(N8471), .A(N8798), .B(N9089));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1969 (.Y(N8739), .A(N8259), .B(N8522));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1970 (.Y(N8586), .A(N8101), .B(N8218));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1971 (.Y(N8317), .A(N8471), .B(N8739));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1972 (.Y(N8432), .A(N8586), .B(N7937));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I1973 (.Y(N8173), .AN(N8870), .B(N8966), .C(N8317), .D(N8668));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1975 (.Y(N7959), .A(N9140), .B(N9004));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1976 (.Y(N8495), .A(N8587), .B(N9034));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1977 (.Y(N7958), .A(N8646), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I10709 (.Y(N8761), .A(N8104), .B(N8035));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1979 (.Y(N8503), .A(N8692), .B(N8770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1980 (.Y(N8070), .A(N7908), .B(N8890));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1981 (.Y(N8338), .A(N8154), .B(N8776));
NAND2X1 inst_cellmath__195__80__2WWMM_2WWMM_I1982 (.Y(N9056), .A(N8166), .B(N8870));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I1983 (.Y(N8886), .A(N9022));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1984 (.Y(N7918), .A(N8886), .B(N7959));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1985 (.Y(N8711), .A(N8070), .B(N8338));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I1986 (.Y(N8562), .A(N8761), .B(N8503), .C(N8495), .D(N7958));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1987 (.Y(N8448), .A(N8001), .B(N8608));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1988 (.Y(N8026), .A(N9056), .B(N8448));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1990 (.Y(N8340), .A(N8931), .B(N9012));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1991 (.Y(N7984), .A(N8043), .B(N9125));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1992 (.Y(N8519), .A(N8795), .B(N9029));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1993 (.Y(N8793), .A(N7978), .B(N9140));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1994 (.Y(N9084), .A(N8927), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1995 (.Y(N8095), .A(N8646), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1996 (.Y(N8357), .A(N8035), .B(N9069));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1997 (.Y(N8618), .A(N8962), .B(N8953));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I1998 (.Y(N8911), .A(N7908), .B(N8187));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I1999 (.Y(N8273), .A(N8970), .B(N8618));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2000 (.Y(N8579), .AN(N8793), .B(N8049), .C(N8001));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2001 (.Y(N8857), .A(N7984), .B(N8048));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2002 (.Y(N7895), .A(N9084), .B(N8095));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2003 (.Y(N8169), .A(N8357), .B(N8519));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2004 (.Y(N8425), .A(N8279), .B(N8911));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2005 (.Y(N8000), .A(N8857), .B(N7895));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2006 (.Y(N8537), .AN(N8340), .B(N8859), .C(N8273));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2007 (.Y(N8123), .A(N8169), .B(N8425));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2008 (.Y(N8638), .A(N8685), .B(N8579), .C(N8000));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2009 (.Y(N8377), .A(N8123), .B(N8537));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2011 (.Y(N8186), .A(N9004), .B(N8205));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2012 (.Y(N8444), .A(N8646), .B(N8178));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2013 (.Y(N9010), .A(N9119), .B(N8854));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2014 (.Y(N8085), .A(N7919), .B(N8274), .C(N8859));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2015 (.Y(N8147), .A(N8912), .B(N8750));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2016 (.Y(N8888), .A(N8724), .B(N8603));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2017 (.Y(N8657), .A(N8186), .B(N8147));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2018 (.Y(N8950), .A(N8281), .B(N9010));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2019 (.Y(N7977), .A(N8362), .B(N8444));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2020 (.Y(N8248), .AN(N8888), .B(N8269), .C(N8550));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2021 (.Y(N8783), .A(N9125), .B(N8795), .C(N8657));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2022 (.Y(N9076), .A(N8950), .B(N7977));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2023 (.Y(N8353), .A(N8085), .B(N8248));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2024 (.Y(N8905), .A(N8783), .B(N9076));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2026 (.Y(N8678), .A(N7911), .B(N8609));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2028 (.Y(N8533), .A(N8837), .B(N8421));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2030 (.Y(N8749), .A(N8678), .B(N8859));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2031 (.Y(N8113), .A(N8603), .B(N9022));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29856 (.Y(N8635), .A(N9109), .B(N9103), .C(N9004), .D(N8646));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2033 (.Y(N8058), .AN(N8530), .B(N8713), .C(N8943));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2034 (.Y(N7962), .A(N8899));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2035 (.Y(N8484), .A(N7962), .B(N8635));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2036 (.Y(N8597), .A(N8749), .B(N8113), .C(N8533));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2037 (.Y(N8325), .A(N8058), .B(N8484));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2039 (.Y(N9035), .A(N8628), .B(N8713));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2040 (.Y(N8652), .A(N9119), .B(N9103));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2041 (.Y(N8194), .A(N8725), .B(N8912));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2042 (.Y(N7968), .A(N8750), .B(N8603));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2043 (.Y(N9067), .A(N8427), .B(N8181), .C(N8481), .D(N8837));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2044 (.Y(N8774), .A(N8652), .B(N7968));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2045 (.Y(N8080), .A(N9067), .B(N8194));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2046 (.Y(N8349), .A(N9035), .B(N8530));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2047 (.Y(N8898), .A(N8646), .B(N8608), .C(N8774));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2048 (.Y(N761), .AN(N8898), .B(N8349), .C(N8080));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2049 (.Y(N8670), .A(N8205), .B(N8116));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2050 (.Y(N8969), .A(N8035), .B(N8943));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2051 (.Y(N8263), .A(N7887), .B(N9119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2052 (.Y(N8712), .A(N8416), .B(N8725));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2053 (.Y(N8802), .A(N8724), .B(N8166));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2054 (.Y(N8106), .A(N8970), .B(N8670));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2055 (.Y(N8624), .A(N8721), .B(N8712));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2056 (.Y(N8920), .A(N8969), .B(N8263));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2057 (.Y(N8478), .AN(N8802), .B(N8837), .C(N8770));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2058 (.Y(N8223), .A(N8106), .B(N8920));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2059 (.Y(N8743), .A(N8478), .B(N8223));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2061 (.Y(N8007), .A(N8713), .B(N8035));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2062 (.Y(N8543), .A(N8481), .B(N8697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2063 (.Y(N8137), .A(N8870), .B(N8572));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2064 (.Y(N8940), .A(N8543), .B(N8620));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2065 (.Y(N7961), .A(N8888), .B(N8523));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2066 (.Y(N8501), .A(N8336));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2067 (.Y(N8407), .A(N8178), .B(N7887), .C(N8501));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2068 (.Y(N8605), .A(N8433), .B(N8407));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2069 (.Y(N9059), .A(N8940), .B(N7961));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2070 (.Y(N8345), .A(N8137), .B(N8007), .C(N9059));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2072 (.Y(N8736), .A(N8608), .B(N8104));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2073 (.Y(N9036), .A(N8943), .B(N8187));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2074 (.Y(N8583), .A(N8550), .B(N8762));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2075 (.Y(N8930), .A(N8859), .B(N8912));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2076 (.Y(N8820), .AN(N8495), .B(N8125), .C(N8659));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2077 (.Y(N8990), .A(N8645), .B(N8583));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2078 (.Y(N8003), .A(N9036), .B(N8685));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2079 (.Y(N8540), .AN(N7940), .B(N8077), .C(N8006));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2081 (.Y(N8380), .A(N8736), .B(N8930));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2083 (.Y(N8094), .A(N8216), .B(N8320), .C(N8380));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2084 (.Y(N8933), .A(N8820), .B(N8094));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2088 (.Y(N8446), .A(N9029), .B(N9052));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2089 (.Y(N8709), .A(N9134), .B(N8646));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2090 (.Y(N9014), .A(N8421), .B(N8953));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2091 (.Y(N8023), .A(N8876), .B(N8481));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2092 (.Y(N8296), .A(N9109), .B(N8947));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2093 (.Y(N8957), .A(N8365), .B(N8446));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29863 (.Y(N7981), .A(N8181), .B(N8049), .C(N7945), .D(N8520));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2095 (.Y(N8516), .A(N8296), .B(N9014), .C(N8023));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2096 (.Y(N8790), .A(N8583), .B(N8712));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2097 (.Y(N9081), .A(N8269), .B(N8457), .C(N8724), .D(N7981));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2098 (.Y(N8089), .A(N8709), .B(N9081));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2099 (.Y(inst_cellmath__197[1]), .A(N8957), .B(N8516), .C(N8790), .D(N8089));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2100 (.Y(N7893), .A(N8043), .B(N8520));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2101 (.Y(N8167), .A(N8001), .B(N8927));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2102 (.Y(N8683), .A(N8427), .B(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2103 (.Y(N8982), .A(N8943), .B(N8692));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2104 (.Y(N8813), .A(N8154), .B(N8603));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2107 (.Y(N8374), .AN(N7990), .B(N9052), .C(N8785));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29864 (.Y(N8636), .A(N8167), .B(N7999), .C(N8683), .D(N7893));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2110 (.Y(N8488), .A(N8813), .B(N8636));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2111 (.Y(N9032), .A(N7887), .B(N8659), .C(N8488));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2114 (.Y(N8016), .A(N8713), .B(N9069));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2115 (.Y(N9130), .A(N8125), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2116 (.Y(N8397), .A(N8697), .B(N8416));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2117 (.Y(N8084), .A(N9022), .B(N9044));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2118 (.Y(N8948), .A(N8962), .B(N9086), .C(N8953), .D(N8876));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2119 (.Y(N7974), .A(N8927), .B(N8274), .C(N9004), .D(N8799));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2120 (.Y(N7930), .A(N8397), .B(N8055));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2121 (.Y(N9073), .A(N8279), .B(N8948));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2122 (.Y(N8461), .A(N8084), .B(N7974));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2123 (.Y(N8903), .A(N9130), .B(N8995), .C(N8016));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2124 (.Y(inst_cellmath__197[3]), .A(N7930), .B(N8903), .C(N9073), .D(N8461));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2125 (.Y(N8974), .A(N8001), .B(N9140));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2126 (.Y(N8805), .A(N8680), .B(N8785));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2127 (.Y(N8460), .A(N8608), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2129 (.Y(N8631), .A(N8207), .B(N8125));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2130 (.Y(N7906), .A(N8659), .B(N8550));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29866 (.Y(N9122), .AN(N8995), .B(N8697), .C(N8460), .D(N8724));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2134 (.Y(N8594), .A(N8185), .B(N8609), .C(N8631));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29865 (.Y(N8872), .A(N7887), .B(N8890), .C(N8776), .D(N8077));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2136 (.Y(N8700), .A(N8805), .B(N8974), .C(N7958));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2139 (.Y(N8390), .AN(N8700), .B(N7906), .C(N7893), .D(N8672));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2142 (.Y(N9064), .A(N8931), .B(N8520));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2143 (.Y(N8458), .A(N8847), .B(N7887));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2144 (.Y(N8719), .A(N9119), .B(N8762));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2145 (.Y(N8414), .AN(N8598), .B(N8104), .C(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2146 (.Y(N8848), .A(N8697), .B(N8870));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2147 (.Y(N8526), .AN(N8090), .B(N8825), .C(N9004));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2148 (.Y(N8669), .A(N8414), .B(N8719));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2149 (.Y(N8968), .A(N8458), .B(N8533));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2150 (.Y(N8262), .A(N8848), .B(N8917), .C(N8741));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2151 (.Y(N8800), .AN(N8859), .B(N9064), .C(N8526));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2152 (.Y(inst_cellmath__197[5]), .A(N8968), .B(N8800), .C(N8262), .D(N8669));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2153 (.Y(N8436), .A(N9012), .B(N8320));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2154 (.Y(N8693), .A(N8608), .B(N8434));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2155 (.Y(N9115), .A(N8365), .B(N8070));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2156 (.Y(N8763), .A(N8436), .B(N9056));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2157 (.Y(N7960), .A(N8188), .B(N8788), .C(N7959), .D(N8645));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2158 (.Y(N8684), .A(N8943), .B(N8953), .C(N8693));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2159 (.Y(N8499), .A(N8816), .B(N8684));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2160 (.Y(inst_cellmath__197[6]), .A(N9115), .B(N7960), .C(N8763), .D(N8499));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2161 (.Y(N7985), .A(N8962), .B(N8481));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2163 (.Y(N8468), .A(N8166), .B(N8603));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2164 (.Y(N9087), .AN(N8572), .B(N8548), .C(N8609));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29867 (.Y(N8733), .AN(N8826), .B(N7908), .C(N8468), .D(N8947));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2166 (.Y(N8619), .A(N8159), .B(N9035));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2167 (.Y(N8213), .A(N7985), .B(N8219), .C(N8668));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2169 (.Y(N8045), .A(N9087), .B(N8619));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2170 (.Y(N8376), .A(N8832), .B(N8659), .C(N8213));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2174 (.Y(N8817), .A(N9034), .B(N8205));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2175 (.Y(N7952), .A(N8363), .B(N9103));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2176 (.Y(N8028), .A(N8724), .B(N8776));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2177 (.Y(N8334), .A(N8962), .B(N7908), .C(N8628), .D(N8035));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2180 (.Y(N7913), .A(N8028), .B(N8631));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29868 (.Y(N8707), .A(N8817), .B(N7952), .C(N7959), .D(N9084));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2182 (.Y(N8022), .A(N8931), .B(N8274), .C(N8859), .D(N7913));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2184 (.Y(N8838), .A(N8362), .B(N8334), .C(N8022));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2187 (.Y(N7890), .A(N8001), .B(N8795));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2191 (.Y(N8907), .A(N8770), .B(N8847));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29869 (.Y(N8726), .A(N8997), .B(N9069), .C(N8457), .D(N8104));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2193 (.Y(N8422), .A(N8544), .B(N8907));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2194 (.Y(N8576), .A(N8912), .B(N8077), .C(N8726));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29870 (.Y(N8855), .A(N9077), .B(N8427), .C(N8799), .D(N8304));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2196 (.Y(N8535), .A(N8697), .B(N8762), .C(N8422));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2197 (.Y(N7998), .A(N8481), .B(N8125), .C(N8855));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2198 (.Y(N8271), .A(N7890), .B(N8793), .C(N8340), .D(N8576));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2201 (.Y(N7947), .A(N7919), .B(N8181));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2204 (.Y(N8329), .A(N8104), .B(N8692));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2205 (.Y(N7910), .A(N9103), .B(N8154));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2206 (.Y(N8702), .A(N8329), .B(N7947));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29871 (.Y(N9126), .A(N8825), .B(N8049), .C(N9125), .D(N9029));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2208 (.Y(N8395), .AN(N7990), .B(N8628), .C(N8178));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2209 (.Y(N8244), .A(N9134), .B(N9034), .C(N8702));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2211 (.Y(N8065), .A(N8659), .B(N7908), .C(N8613));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2212 (.Y(N7970), .A(N8802), .B(N8065));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2214 (.Y(N9009), .A(N8603), .B(N9044), .C(N7970));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2215 (.Y(N8779), .A(N8395), .B(N9009));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2217 (.Y(N8204), .A(N8653), .B(N7919));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2218 (.Y(N8723), .A(N8520), .B(N8997));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2219 (.Y(N9025), .A(N9029), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2220 (.Y(N7886), .A(N9119), .B(N8187));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2221 (.Y(N8675), .A(N9071), .B(N8204));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2222 (.Y(N8971), .A(N8762), .B(N8725));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2223 (.Y(N8922), .AN(N8964), .B(N8962), .C(N8692));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2224 (.Y(N9097), .A(N8917), .B(N7886));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2225 (.Y(N8627), .A(N9025), .B(N7933));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2226 (.Y(N7941), .A(N8922), .B(N8971));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2227 (.Y(N8479), .A(N8116), .B(N8587), .C(N8870), .D(N9097));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2229 (.Y(N8319), .AN(N7941), .B(N8340), .C(N8761), .D(N8723));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2232 (.Y(N8998), .A(N7919), .B(N8520));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2233 (.Y(N8008), .A(N8001), .B(N7945));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2234 (.Y(N8283), .A(N9029), .B(N9034));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2235 (.Y(N8827), .A(N8876), .B(N7887));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2237 (.Y(N8388), .A(N8659), .B(N9103));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29872 (.Y(N9062), .A(N8890), .B(N8725), .C(N8697), .D(N9119));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2242 (.Y(N8075), .A(N8283), .B(N8827));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2243 (.Y(N8346), .AN(N9130), .B(N8912), .C(N9022));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29873 (.Y(N8455), .A(N8008), .B(N8388), .C(N8998), .D(N8503));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2245 (.Y(N8895), .A(N9062), .B(N8075));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2249 (.Y(N8413), .A(N8520), .B(N7945));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2250 (.Y(N7988), .A(N8205), .B(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2251 (.Y(N8260), .A(N8116), .B(N8320));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2252 (.Y(N8102), .A(N7908), .B(N8854));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2253 (.Y(N8360), .A(N8207), .B(N8724));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2254 (.Y(N9008), .A(N8572), .B(N8109));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2255 (.Y(N8472), .A(N8793), .B(N8413), .C(N7988), .D(N8532));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2258 (.Y(N8316), .A(N8491), .B(N8260));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2259 (.Y(N8174), .A(N9008), .B(N8472));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29875 (.Y(N8864), .A(N8982), .B(N8360), .C(N8102), .D(N8706));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2261 (.Y(N8655), .A(N8316), .B(N9022), .C(N8776));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2265 (.Y(N8383), .A(N9092), .B(N8043));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2266 (.Y(N8644), .A(N8049), .B(N8997));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2267 (.Y(N7957), .A(N9140), .B(N8097));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2268 (.Y(N8494), .A(N8066), .B(N8104));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2269 (.Y(N8887), .AN(N8598), .B(N8659), .C(N8890));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2272 (.Y(N8960), .AN(N8494), .B(N8201), .C(N8854));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2273 (.Y(N9138), .AN(N8712), .B(N9109), .C(N8750), .D(N8569));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29876 (.Y(N8153), .A(N8644), .B(N8008), .C(N7957), .D(N8132));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2275 (.Y(N7983), .A(N8960), .B(N8153));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2276 (.Y(N9085), .AN(N8859), .B(N8383), .C(N9138));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2277 (.Y(N8352), .A(N8269), .B(N9012), .C(N7983));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2280 (.Y(N8042), .A(N8274), .B(N8997));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2281 (.Y(N8858), .A(N8178), .B(N8962));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2282 (.Y(N8611), .A(N8770), .B(N7887));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2283 (.Y(N8986), .A(N8753), .B(N8042));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2284 (.Y(N8538), .A(N9140), .B(N8927), .C(N8077));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2285 (.Y(N8815), .A(N8858), .B(N7886));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2286 (.Y(N8124), .AN(N8538), .B(N8205), .C(N8035));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2288 (.Y(N7950), .A(N8611), .B(N7933), .C(N8930));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2292 (.Y(N8952), .A(N8628), .B(N8943));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2294 (.Y(N8835), .A(N9119), .B(N8659));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2295 (.Y(N8951), .A(N8859), .B(N8416));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2296 (.Y(N8400), .A(N8870), .B(N8109));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2297 (.Y(N8656), .A(N9140), .B(N8725), .C(N8825), .D(N8724));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2298 (.Y(N8086), .A(N8952), .B(N8656));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29877 (.Y(N8784), .A(N8421), .B(N8320), .C(N8205), .D(N7887));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2300 (.Y(N8514), .A(N8400), .B(N8835));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2301 (.Y(inst_cellmath__197[16]), .A(N8951), .B(N8784), .C(N8514), .D(N8086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2302 (.Y(N8307), .A(N8205), .B(N8427));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2303 (.Y(N9043), .A(N8628), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2304 (.Y(N8165), .A(N8770), .B(N8481));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2305 (.Y(N8980), .A(N8750), .B(N8724));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2306 (.Y(N8563), .A(N9022), .B(N8572));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2307 (.Y(N8714), .A(N8077), .B(N8109));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2308 (.Y(N8808), .A(N8307), .B(N8615));
INVXL inst_cellmath__195__80__2WWMM_2WWMM_I2311 (.Y(N8371), .A(N8165));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29878 (.Y(N8326), .A(N8969), .B(N8824), .C(N8563), .D(N8194));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29879 (.Y(N8596), .AN(N8714), .B(N8980), .C(N8326), .D(N9043));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2315 (.Y(N8485), .AN(N8835), .B(N8304), .C(N8608));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2320 (.Y(N8549), .A(N8304), .B(N8646));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2321 (.Y(N8775), .AN(N8549), .B(N7919), .C(N8205));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2322 (.Y(N7926), .AN(N8980), .B(N8077), .C(N8572));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2323 (.Y(N8081), .A(N8712), .B(N8824));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2324 (.Y(N8720), .A(N8460), .B(N8081));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2325 (.Y(N8034), .A(N8969), .B(N8611), .C(N8113), .D(N8775));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2328 (.Y(N9095), .A(N8178), .B(N8837));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2329 (.Y(N8477), .A(N9095), .B(N8620));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2330 (.Y(N9042), .A(N8007), .B(N8523));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2331 (.Y(N8052), .A(N8888), .B(N8137));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2332 (.Y(N8589), .A(N8953), .B(N7887), .C(N8477));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2333 (.Y(N8695), .AN(N8501), .B(N8543), .C(N8433));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2338 (.Y(N8717), .A(N8799), .B(N8304));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29880 (.Y(N8453), .A(N9077), .B(N8825), .C(N8434), .D(N8181));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2341 (.Y(N8303), .A(N9029), .B(N9140), .C(N8453));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2342 (.Y(N8566), .A(N8563), .B(N8888));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2343 (.Y(N8843), .A(N8441), .B(N8309), .C(N8523), .D(N8717));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2344 (.Y(N8157), .A(N8011), .B(N8296), .C(N8021));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2345 (.Y(N8410), .A(N8303), .B(N9104));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2346 (.Y(inst_cellmath__195[0]), .A(N8157), .B(N8843), .C(N8410), .D(N8566));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2347 (.Y(N8313), .A(N7887), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2348 (.Y(N7899), .A(N8724), .B(N9022));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2349 (.Y(N8689), .A(N8672), .B(N7882));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2350 (.Y(N8991), .A(N8927), .B(N9140), .C(N9134), .D(N9125));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2351 (.Y(N8002), .A(N8545), .B(N8077));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2352 (.Y(N8277), .AN(N8309), .B(N8456), .C(N8002));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2353 (.Y(N8819), .A(N8697), .B(N8363), .C(N8689));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2354 (.Y(N8935), .AN(N9020), .B(N8097), .C(N8628));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2355 (.Y(N8379), .A(N8130), .B(N8991));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2356 (.Y(N8492), .A(N7899), .B(N8159));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2357 (.Y(N7953), .A(N8935), .B(N8313));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2358 (.Y(N8234), .A(N8277), .B(N8819));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2359 (.Y(inst_cellmath__195[1]), .A(N8379), .B(N8492), .C(N7953), .D(N8234));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2360 (.Y(N8297), .A(N8795), .B(N8799));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2361 (.Y(N8150), .A(N8947), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2362 (.Y(N9139), .A(N8762), .B(N8154));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2363 (.Y(N8663), .A(N8309), .B(N8150));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2364 (.Y(N8789), .A(N7947), .B(N8297));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2365 (.Y(N8091), .A(N9052), .B(N9034), .C(N8663));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2366 (.Y(N8616), .A(N8002), .B(N8789));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2367 (.Y(N9030), .AN(N8712), .B(N8750), .C(N8870));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2368 (.Y(N8727), .A(N8616), .B(N8270), .C(N9139));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2370 (.Y(N8038), .A(N8320), .B(N8770), .C(N8727));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2373 (.Y(N8812), .A(N9034), .B(N8304));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2375 (.Y(N7898), .A(N8953), .B(N8569));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2376 (.Y(N8331), .AN(N8309), .B(N8947), .C(N8832));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2377 (.Y(N8063), .AN(N7898), .B(N7945), .C(N8795));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2381 (.Y(N8442), .A(N8362), .B(N8209));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29883 (.Y(N8290), .AN(N8331), .B(N8178), .C(N8442), .D(N8066));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2379 (.Y(N8879), .A(N8812), .B(N7959));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2380 (.Y(N8184), .A(N8194), .B(N8063));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2382 (.Y(N8017), .A(N9008), .B(N8879));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2384 (.Y(N8978), .A(N7908), .B(N9119), .C(N8184));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2388 (.Y(N9074), .A(N8653), .B(N9092));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2389 (.Y(N7929), .A(N8104), .B(N8876));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2390 (.Y(N9027), .A(N9109), .B(N8832));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2391 (.Y(N8852), .A(N8365), .B(N7893));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2392 (.Y(N8163), .A(N8463), .B(N8777), .C(N9074));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2393 (.Y(N8418), .A(N7929), .B(N8934));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2394 (.Y(N8976), .A(N9052), .B(N8097), .C(N8418));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2395 (.Y(N8266), .A(N8002), .B(N8163));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2397 (.Y(N8634), .A(N9027), .B(N8603), .C(N8852));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2400 (.Y(N8322), .A(N8653), .B(N8043));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2401 (.Y(N8593), .A(N9134), .B(N8587));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2402 (.Y(N8874), .A(N8320), .B(N8713));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2403 (.Y(N8180), .A(N8434), .B(N8943));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2404 (.Y(N8699), .A(N8890), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2405 (.Y(N9002), .A(N8659), .B(N8750));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29884 (.Y(N9121), .A(N8309), .B(N8593), .C(N8699), .D(N8322));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2414 (.Y(N9024), .A(N9069), .B(N8943));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2415 (.Y(N8527), .A(N8837), .B(N9086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2416 (.Y(N8408), .A(N8953), .B(N8770));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2417 (.Y(N8364), .A(N8408), .B(N8188));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2418 (.Y(N8221), .A(N8467), .B(N8527), .C(N8683));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2421 (.Y(N8051), .A(N7945), .B(N8587), .C(N8035), .D(N8364));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29885 (.Y(N7938), .A(N8095), .B(N8279), .C(N9024), .D(N8117));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29886 (.Y(N8318), .AN(N8221), .B(N9056), .C(N8051), .D(N8563));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2425 (.Y(N9041), .A(N8998), .B(N8365), .C(N7938));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2427 (.Y(inst_cellmath__195[6]), .A(N9041), .B(N8318));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2428 (.Y(N8005), .A(N8927), .B(N8039));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2429 (.Y(N9116), .A(N9069), .B(N8962));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2430 (.Y(N8745), .A(N8187), .B(N8207));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2431 (.Y(N8237), .A(N8166), .B(N9022));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2432 (.Y(N8498), .A(N9116), .B(N8949));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2435 (.Y(N8343), .A(N8569), .B(N7908), .C(N8498));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2436 (.Y(N8604), .AN(N8408), .B(N8116), .C(N8178));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29887 (.Y(N8893), .A(N8593), .B(N7988), .C(N8745), .D(N8005));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2438 (.Y(N8451), .A(N8237), .B(N8893));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2440 (.Y(N8324), .A(N8363), .B(N8762), .C(N8451));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29888 (.Y(inst_cellmath__195[7]), .A(N8343), .B(N8604), .C(N8930), .D(N8324));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2443 (.Y(N8098), .A(N8288), .B(N8609));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2444 (.Y(N8621), .A(N8628), .B(N9069));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2445 (.Y(N8734), .A(N9103), .B(N8603));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2446 (.Y(N8860), .A(N8181), .B(N7978), .C(N8098));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2447 (.Y(N8171), .AN(N7898), .B(N8587), .C(N9027), .D(N8039));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2450 (.Y(N8012), .A(N7962), .B(N8104), .C(N8837));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2451 (.Y(N8127), .A(N8911), .B(N8012));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29889 (.Y(N8539), .A(N8734), .B(N8621), .C(N8860), .D(N8171));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2453 (.Y(N9110), .A(N8383), .B(N8365), .C(N8539));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2454 (.Y(inst_cellmath__195[8]), .A(N8127), .B(N9110));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2455 (.Y(N8335), .A(N7919), .B(N9125));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2457 (.Y(N7914), .A(N8785), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2459 (.Y(N8708), .A(N8201), .B(N8481));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2460 (.Y(N8403), .AN(N8335), .B(N8997), .C(N9029));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2461 (.Y(N8294), .A(N8859), .B(N8166));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29890 (.Y(N8955), .A(N8587), .B(N9086), .C(N9052), .D(N8104));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2465 (.Y(N7980), .A(N8955), .B(N7910));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29891 (.Y(N8250), .A(N8721), .B(N7914), .C(N8708), .D(N8403));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29892 (.Y(inst_cellmath__195[9]), .A(N8294), .B(N8606), .C(N7980), .D(N8250));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2472 (.Y(N9105), .A(N8001), .B(N9029), .C(N8077));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29893 (.Y(N8373), .A(N8205), .B(N8434), .C(N9109), .D(N8207));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2475 (.Y(N9048), .AN(N8028), .B(N8770), .C(N7908));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29894 (.Y(N8061), .AN(N8373), .B(N9014), .C(N9048), .D(N8995));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2477 (.Y(N8752), .A(N9139), .B(N9105));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2479 (.Y(N8328), .AN(N8752), .B(N8928), .C(N8495), .D(N8609));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2480 (.Y(inst_cellmath__195[10]), .A(N8061), .B(N8328));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2481 (.Y(N8302), .A(N8799), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2482 (.Y(N8552), .A(N8205), .B(N8628));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2483 (.Y(N8144), .A(N8837), .B(N8962));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2484 (.Y(N8394), .A(N8421), .B(N9086));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2485 (.Y(N8778), .A(N8187), .B(N8832));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2486 (.Y(N8245), .A(N8274), .B(N8692), .C(N9077), .D(N9125));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2487 (.Y(N8350), .A(N8394), .B(N8302));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2488 (.Y(N7927), .A(N8778), .B(N8245));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2489 (.Y(N8082), .A(N8967), .B(N8552));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2490 (.Y(N8614), .A(N8350), .B(N8144));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2491 (.Y(N8900), .A(N8270), .B(N8829));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2492 (.Y(inst_cellmath__195[11]), .A(N8614), .B(N8900), .C(N8082), .D(N7927));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2493 (.Y(N8674), .A(N8680), .B(N8608));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2494 (.Y(N9098), .A(N8653), .B(N9119));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2495 (.Y(N8480), .AN(N8329), .B(N9029), .C(N8799));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2496 (.Y(N9045), .A(N8745), .B(N8672), .C(N8219));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2499 (.Y(N8009), .A(N8870), .B(N8077), .C(N9045));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2500 (.Y(N8696), .A(N8055), .B(N8527), .C(N8480), .D(N9043));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29896 (.Y(N8999), .A(N8674), .B(N9139), .C(N7906), .D(N9098));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2502 (.Y(N8282), .A(N8009), .B(N8999));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2503 (.Y(inst_cellmath__195[12]), .A(N8696), .B(N8282));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2504 (.Y(N8505), .A(N8795), .B(N7978));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2505 (.Y(N8160), .A(N7908), .B(N9103));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2506 (.Y(N9023), .A(N8672), .B(N8335));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2507 (.Y(N8568), .A(N9080), .B(N8505));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2508 (.Y(N7883), .A(N8692), .B(N8481), .C(N8724), .D(N8154));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2509 (.Y(N8524), .A(N7976), .B(N7971), .C(N8160), .D(N8939));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2510 (.Y(N9090), .A(N8603), .B(N8870), .C(N8460));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2511 (.Y(N8946), .A(N8524), .B(N8568), .C(N9023));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2512 (.Y(N8361), .A(N8357), .B(N8946));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2513 (.Y(N8103), .A(N7883), .B(N8563), .C(N9090));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2514 (.Y(inst_cellmath__195[13]), .A(N8361), .B(N8103));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2515 (.Y(N8473), .A(N8043), .B(N8049));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2517 (.Y(N7901), .A(N8434), .B(N8876));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2518 (.Y(N8772), .A(N8187), .B(N9109));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29897 (.Y(N8938), .AN(N9071), .B(N8997), .C(N8643), .D(N7945));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2520 (.Y(N8823), .A(N8365), .B(N7901));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2521 (.Y(N9113), .A(N8473), .B(N8505));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2522 (.Y(N8133), .A(N8386), .B(N8647));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2523 (.Y(N8384), .A(N7959), .B(N8772));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2525 (.Y(N8496), .A(N8166), .B(N8077), .C(N8384));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2526 (.Y(N8071), .AN(N8162), .B(N8097), .C(N8035));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2528 (.Y(N8610), .A(N9113), .B(N8133), .C(N8823));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29898 (.Y(inst_cellmath__195[14]), .A(N8938), .B(N8071), .C(N8496), .D(N8610));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2531 (.Y(N8029), .A(N9004), .B(N8039));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2532 (.Y(N8841), .A(N8178), .B(N9077));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2533 (.Y(N8254), .A(N8166), .B(N8572));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2534 (.Y(N8730), .A(N8077), .B(N9044));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2535 (.Y(N8794), .AN(N8042), .B(N8269), .C(N8653));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2536 (.Y(N8212), .A(N8732), .B(N8029), .C(N7997));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2537 (.Y(N9033), .A(N8801), .B(N8147), .C(N8730));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2538 (.Y(N7896), .A(N8096), .B(N8794), .C(N8254));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2539 (.Y(N8580), .A(N8517), .B(N8841), .C(N8966));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2540 (.Y(N8305), .A(N8953), .B(N8481), .C(N8212));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2541 (.Y(N8426), .A(N8028), .B(N8305));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2542 (.Y(inst_cellmath__195[15]), .A(N9033), .B(N8580), .C(N7896), .D(N8426));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2543 (.Y(N8639), .A(N9092), .B(N8997));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2544 (.Y(N8232), .A(N9052), .B(N8680));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2545 (.Y(N8242), .A(N8304), .B(N8456));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2546 (.Y(N9051), .A(N8943), .B(N8421));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2547 (.Y(N8881), .A(N8598), .B(N8639));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2548 (.Y(N9133), .A(N8725), .B(N8216));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2549 (.Y(N8292), .AN(N8242), .B(N7978), .C(N8927));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2551 (.Y(N8401), .AN(N8817), .B(N8187), .C(N8890));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2552 (.Y(N8555), .A(N8292), .B(N9051));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29903 (.Y(N8658), .AN(N8881), .B(N7890), .C(N8401), .D(N8232));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2554 (.Y(N8148), .A(N9133), .B(N8458));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2556 (.Y(inst_cellmath__195[16]), .A(N8951), .B(N8148), .C(N8555), .D(N8658));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2557 (.Y(N8308), .A(N8890), .B(N8207));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2558 (.Y(N8679), .A(N8947), .B(N8962), .C(N8457), .D(N8653));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2559 (.Y(N7996), .A(N8132), .B(N7948));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2560 (.Y(N8268), .A(N8433), .B(N8362));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2561 (.Y(N9102), .A(N9056), .B(N8276));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2562 (.Y(N8114), .A(N7996), .B(N8268));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2563 (.Y(N8372), .A(N8308), .B(N8679), .C(N8534), .D(N8114));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2564 (.Y(inst_cellmath__195[17]), .A(N9102), .B(N8372));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2565 (.Y(N8064), .A(N8832), .B(N8363));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2566 (.Y(N8013), .A(N8859), .B(N8750));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2567 (.Y(N9124), .A(N8394), .B(N8064));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2568 (.Y(N8393), .A(N8142), .B(N9124));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2569 (.Y(N7993), .A(N8825), .B(N9029), .C(N8393));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2570 (.Y(N8243), .A(N8721), .B(N7993));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2571 (.Y(N8508), .A(N8758), .B(N8007));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2572 (.Y(N9068), .A(N8013), .B(N8028), .C(N8165));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2573 (.Y(N8612), .A(N8753), .B(N7997), .C(N8260), .D(N9064));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2574 (.Y(inst_cellmath__195[18]), .A(N8508), .B(N9068), .C(N8612), .D(N8243));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2575 (.Y(N8571), .A(N9029), .B(N9134));
AND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2576 (.Y(N7884), .A(N8785), .B(N8205));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2577 (.Y(N8671), .A(N8931), .B(N8035));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2578 (.Y(N8528), .A(N8876), .B(N9109));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2579 (.Y(N8107), .A(N8859), .B(N8724));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2580 (.Y(N8625), .A(N8886), .B(N8494));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2581 (.Y(N8921), .A(N8528), .B(N8571));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2582 (.Y(N8744), .A(N8947), .B(N8207), .C(N8921));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I2583 (.Y(N8053), .AN(N9043), .B(N8692), .C(N7884), .D(N8421));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2584 (.Y(N8590), .A(N8495), .B(N8408), .C(N9139));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2585 (.Y(N8867), .A(N8671), .B(N8744));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2586 (.Y(N7903), .A(N8053), .B(N8107));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2587 (.Y(inst_cellmath__195[19]), .A(N8625), .B(N8867), .C(N7903), .D(N8590));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2588 (.Y(N8138), .A(N8457), .B(N7919));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2589 (.Y(N8502), .A(N8628), .B(N8434));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2590 (.Y(N8767), .A(N9077), .B(N8953));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2591 (.Y(N8074), .A(N8481), .B(N8854));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2594 (.Y(N8454), .A(N8048), .B(N8233));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29906 (.Y(N8844), .A(N8777), .B(N8928), .C(N8138), .D(N8767));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2598 (.Y(N9142), .A(N8502), .B(N8074));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2599 (.Y(N8158), .A(N8370), .B(N8441), .C(N9020), .D(N8844));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29908 (.Y(N8411), .A(N8776), .B(N8109), .C(N8302), .D(N8454));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2601 (.Y(inst_cellmath__195[20]), .A(N7909), .B(N9142), .C(N8158), .D(N8411));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2602 (.Y(N8584), .A(N8125), .B(N8550));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2603 (.Y(N8992), .A(N8970), .B(N8584));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2604 (.Y(N9111), .AN(N7990), .B(N9052), .C(N8795));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2605 (.Y(N8936), .A(N8901), .B(N8598), .C(N9091));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2606 (.Y(N8821), .A(N8533), .B(N8028));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2609 (.Y(N8919), .A(N8481), .B(N9119), .C(N7909));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2610 (.Y(N9053), .A(N9111), .B(N8919));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29910 (.Y(N8759), .A(N8936), .B(N8992), .C(N7962), .D(N8821));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2612 (.Y(inst_cellmath__195[21]), .A(N9053), .B(N8759));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2613 (.Y(N8192), .A(N8520), .B(N8001));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2614 (.Y(N8024), .A(N8608), .B(N8178));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2615 (.Y(N8151), .A(N8154), .B(N8697));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2616 (.Y(N8405), .A(N8416), .B(N8724));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2617 (.Y(N8662), .A(N8776), .B(N8603));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2618 (.Y(N8958), .A(N8545), .B(N9044));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2619 (.Y(N8252), .A(N8392), .B(N8192));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2620 (.Y(N8909), .A(N8252), .B(N7884));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2623 (.Y(N8040), .A(N8549), .B(N8283), .C(N8611));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2624 (.Y(N7934), .A(N8909), .B(N8662));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2625 (.Y(N8210), .A(N8405), .B(N8527));
OR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I29913 (.Y(N8465), .A(N8958), .B(N8151), .C(N8764), .D(N8102));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2627 (.Y(N8728), .A(N8024), .B(N8465));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2628 (.Y(inst_cellmath__195[22]), .A(N8210), .B(N8040), .C(N7934), .D(N8728));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2632 (.Y(N8121), .A(N8876), .B(N8569));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29914 (.Y(N8489), .A(N8181), .B(N7978), .C(N7945), .D(N8201));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2635 (.Y(N8755), .A(N8723), .B(N8121));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2636 (.Y(N8183), .A(N8116), .B(N8890), .C(N8854), .D(N8304));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2638 (.Y(N8880), .A(N9140), .B(N8799), .C(N8755));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2639 (.Y(N9007), .AN(N8958), .B(N8587), .C(N8680));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29915 (.Y(N8704), .A(N8697), .B(N8912), .C(N8064), .D(N8489));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29916 (.Y(N8553), .AN(N8183), .B(N8178), .C(N8704), .D(N8434));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2642 (.Y(N8018), .A(N9007), .B(N8362));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2643 (.Y(N8834), .AN(N8880), .B(N8776), .C(N8870));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2645 (.Y(N9131), .A(N8834), .B(N8553));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2646 (.Y(inst_cellmath__195[23]), .A(N8018), .B(N9131));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2648 (.Y(N8531), .AN(N8598), .B(N8049), .C(N7978));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2649 (.Y(N8924), .A(N8274), .B(N8825), .C(N8859));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2651 (.Y(N8975), .A(N8812), .B(N8308));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2653 (.Y(N8369), .AN(N8975), .B(N8441), .C(N8340), .D(N7952));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29918 (.Y(N8632), .AN(N8886), .B(N7919), .C(N8369), .D(N9092));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2652 (.Y(N8267), .A(N8772), .B(N8029), .C(N8408));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2656 (.Y(N8747), .A(N8924), .B(N8028), .C(N8531));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29919 (.Y(inst_cellmath__195[24]), .AN(N8632), .B(N8693), .C(N8747), .D(N8267));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2659 (.Y(N8348), .A(N8572), .B(N9044));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2660 (.Y(N8650), .A(N8825), .B(N8520), .C(N8626));
NAND3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2661 (.Y(N7966), .AN(N8974), .B(N9086), .C(N8953));
NOR3XL inst_cellmath__195__80__2WWMM_2WWMM_I2662 (.Y(N9065), .A(N8772), .B(N8995), .C(N8096));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2663 (.Y(N8588), .A(N8770), .B(N8207), .C(N8569));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2664 (.Y(N8079), .A(N8227), .B(N8588));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2665 (.Y(N8459), .A(N8348), .B(N7966));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2666 (.Y(N8897), .A(N8113), .B(N8824));
NOR3BXL inst_cellmath__195__80__2WWMM_2WWMM_I2667 (.Y(N7925), .AN(N9065), .B(N8242), .C(N8650));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2668 (.Y(inst_cellmath__195[25]), .A(N8079), .B(N8459), .C(N7925), .D(N8897));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2670 (.Y(N8222), .A(N8997), .B(N9092), .C(N8520), .D(N8304));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29920 (.Y(N8050), .AN(N9002), .B(N8847), .C(N8501), .D(N8178));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29921 (.Y(N8176), .AN(N8460), .B(N8222), .C(N8050), .D(N8631));
NOR4X1 inst_cellmath__195__80__2WWMM_2WWMM_I2675 (.Y(N8437), .A(N7886), .B(N8816), .C(N8491), .D(N8662));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2677 (.Y(inst_cellmath__195[26]), .A(N8437), .B(N8176));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2678 (.Y(N7920), .A(N8943), .B(N8770));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2680 (.Y(N8892), .A(N9091), .B(N8841));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29922 (.Y(N8565), .AN(N9056), .B(N7887), .C(N7962), .D(N8187));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2683 (.Y(N8031), .A(N7940), .B(N8563));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2685 (.Y(N8409), .AN(N8031), .B(N7911), .C(N7920), .D(N8717));
NAND4BXL inst_cellmath__195__80__2WWMM_2WWMM_I29924 (.Y(inst_cellmath__195[27]), .AN(N8565), .B(N8714), .C(N8409), .D(N8892));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2688 (.Y(N8913), .A(N8456), .B(N8066));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2689 (.Y(N8215), .A(N8770), .B(N9119));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2690 (.Y(N8046), .A(N9022), .B(N8545));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2691 (.Y(N8582), .A(N7911), .B(N8549));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2692 (.Y(N8687), .A(N8712), .B(N8913));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2695 (.Y(N8128), .A(N7940), .B(N8046));
AND4XL inst_cellmath__195__80__2WWMM_2WWMM_I29926 (.Y(N8640), .A(N8468), .B(N8714), .C(N8582), .D(N8687));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I2697 (.Y(N8378), .AN(N8128), .B(N8276), .C(N8215), .D(N8362));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2698 (.Y(inst_cellmath__195[28]), .A(N8640), .B(N8378));
NAND2XL inst_cellmath__195__80__2WWMM_2WWMM_I2699 (.Y(N8067), .A(N8795), .B(N8304));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2701 (.Y(N8839), .A(N8132), .B(N8730));
NAND3XL inst_cellmath__195__80__2WWMM_2WWMM_I2704 (.Y(N8956), .A(N8697), .B(N9119), .C(N8839));
NOR4BX1 inst_cellmath__195__80__2WWMM_2WWMM_I29928 (.Y(N8786), .AN(N8371), .B(N8194), .C(N8956), .D(N8067));
NOR2XL inst_cellmath__195__80__2WWMM_2WWMM_I2703 (.Y(N8404), .A(N8362), .B(N9056));
NAND4XL inst_cellmath__195__80__2WWMM_2WWMM_I2706 (.Y(inst_cellmath__195[29]), .A(N8128), .B(N8404), .C(N7962), .D(N8786));
INVX3 inst_cellmath__198_0_I2708 (.Y(N10418), .A(inst_cellmath__61[1]));
CLKINVX12 inst_cellmath__198_0_I2711 (.Y(N10622), .A(inst_cellmath__61[2]));
INVX3 inst_cellmath__198_0_I2713 (.Y(N10810), .A(inst_cellmath__61[3]));
INVX3 inst_cellmath__198_0_I2714 (.Y(N10867), .A(inst_cellmath__61[4]));
INVX3 inst_cellmath__198_0_I2715 (.Y(N10431), .A(inst_cellmath__61[5]));
CLKINVX6 inst_cellmath__198_0_I2720 (.Y(N10634), .A(N3808));
INVX2 inst_cellmath__198_0_I2724 (.Y(N10823), .A(inst_cellmath__61[7]));
INVX1 inst_cellmath__198_0_I29260 (.Y(N44729), .A(N10823));
INVX2 inst_cellmath__198_0_I29261 (.Y(N44730), .A(N44729));
INVX3 inst_cellmath__198_0_I2728 (.Y(N11027), .A(inst_cellmath__61[8]));
INVX3 inst_cellmath__198_0_I2730 (.Y(N10590), .A(inst_cellmath__61[9]));
INVX2 inst_cellmath__198_0_I2735 (.Y(N10542), .A(inst_cellmath__61[12]));
INVX2 inst_cellmath__198_0_I2736 (.Y(N10727), .A(inst_cellmath__61[13]));
INVX3 inst_cellmath__198_0_I2737 (.Y(N10922), .A(inst_cellmath__61[14]));
INVX3 inst_cellmath__198_0_I2739 (.Y(N10491), .A(inst_cellmath__61[15]));
INVX3 inst_cellmath__198_0_I2741 (.Y(N10551), .A(inst_cellmath__115__W1[0]));
INVX3 inst_cellmath__198_0_I2743 (.Y(N10878), .A(inst_cellmath__61[0]));
NOR2XL inst_cellmath__198_0_I2750 (.Y(N10481), .A(N10878), .B(N10810));
NOR2XL inst_cellmath__198_0_I2751 (.Y(N10749), .A(N10878), .B(N10867));
NOR2XL inst_cellmath__198_0_I2752 (.Y(N11037), .A(N10878), .B(N10431));
NOR2XL inst_cellmath__198_0_I2753 (.Y(N10676), .A(N10878), .B(N10634));
NOR2XL inst_cellmath__198_0_I2754 (.Y(N10947), .A(N10878), .B(N44730));
NOR2XL inst_cellmath__198_0_I2755 (.Y(N10600), .A(N10878), .B(N11027));
NOR2XL inst_cellmath__198_0_I2756 (.Y(N10865), .A(N10878), .B(N10590));
NOR2XL inst_cellmath__198_0_I2757 (.Y(N10516), .A(N10878), .B(N3809));
NOR2XL inst_cellmath__198_0_I2758 (.Y(N10781), .A(N10878), .B(N10973));
NOR2XL inst_cellmath__198_0_I2759 (.Y(N10428), .A(N10878), .B(N10542));
NOR2XL inst_cellmath__198_0_I2760 (.Y(N10706), .A(N10878), .B(N10727));
NOR2XL inst_cellmath__198_0_I2761 (.Y(N10987), .A(N10878), .B(N10922));
NOR2X2 inst_cellmath__198_0_I2762 (.Y(N10630), .A(N10878), .B(N10491));
OR2XL inst_cellmath__198_0_I2763 (.Y(N10673), .A(N10878), .B(N10551));
NOR2XL inst_cellmath__198_0_I2764 (.Y(N10587), .A(N10622), .B(N10418));
NOR2XL inst_cellmath__198_0_I2765 (.Y(N10852), .A(N10418), .B(N10810));
NOR2XL inst_cellmath__198_0_I2766 (.Y(N10504), .A(N10418), .B(N10867));
NOR2XL inst_cellmath__198_0_I2767 (.Y(N10765), .A(N10431), .B(N10418));
NOR2XL inst_cellmath__198_0_I2768 (.Y(N10415), .A(N10634), .B(N10418));
NOR2XL inst_cellmath__198_0_I2769 (.Y(N10693), .A(N10418), .B(N44730));
NOR2XL inst_cellmath__198_0_I2770 (.Y(N10970), .A(N10418), .B(N11027));
NOR2XL inst_cellmath__198_0_I2771 (.Y(N10619), .A(N10418), .B(N10590));
NOR2XL inst_cellmath__198_0_I2772 (.Y(N10889), .A(N3809), .B(N10418));
NOR2XL inst_cellmath__198_0_I2773 (.Y(N10538), .A(N10418), .B(N10973));
NOR2XL inst_cellmath__198_0_I2774 (.Y(N10804), .A(N10418), .B(N10542));
NOR2XL inst_cellmath__198_0_I2775 (.Y(N10451), .A(N10727), .B(N10418));
NOR2XL inst_cellmath__198_0_I2776 (.Y(N10722), .A(N10922), .B(N10418));
NOR2XL inst_cellmath__198_0_I2777 (.Y(N11007), .A(N10491), .B(N10418));
OR2XL inst_cellmath__198_0_I11210 (.Y(N10805), .A(N10551), .B(N10418));
NOR2XL inst_cellmath__198_0_I2779 (.Y(N10953), .A(N10622), .B(N10810));
NOR2XL inst_cellmath__198_0_I2780 (.Y(N10605), .A(N10622), .B(N10867));
NOR2XL inst_cellmath__198_0_I2781 (.Y(N10874), .A(N10622), .B(N10431));
NOR2XL inst_cellmath__198_0_I2782 (.Y(N10523), .A(N10622), .B(N10634));
NOR2XL inst_cellmath__198_0_I2783 (.Y(N10788), .A(N10622), .B(N44730));
NOR2XL inst_cellmath__198_0_I2784 (.Y(N10436), .A(N10622), .B(N11027));
NOR2XL inst_cellmath__198_0_I2785 (.Y(N10712), .A(N10622), .B(N10590));
NOR2XL inst_cellmath__198_0_I2786 (.Y(N10994), .A(N10622), .B(N3809));
NOR2XL inst_cellmath__198_0_I2787 (.Y(N10637), .A(N10622), .B(N10973));
NOR2XL inst_cellmath__198_0_I2788 (.Y(N10907), .A(N10622), .B(N10542));
NOR2XL inst_cellmath__198_0_I2789 (.Y(N10560), .A(N10622), .B(N10727));
NOR2XL inst_cellmath__198_0_I2790 (.Y(N10827), .A(N10622), .B(N10922));
NOR2XL inst_cellmath__198_0_I2791 (.Y(N10476), .A(N10622), .B(N10491));
OR2XL inst_cellmath__198_0_I2792 (.Y(N10944), .A(N10622), .B(N10551));
INVXL inst_cellmath__198_0_I2793 (.Y(N10510), .A(N10810));
NOR2XL inst_cellmath__198_0_I2794 (.Y(N10422), .A(N10867), .B(N10810));
NOR2XL inst_cellmath__198_0_I2795 (.Y(N10699), .A(N10810), .B(N10431));
NOR2XL inst_cellmath__198_0_I2796 (.Y(N10979), .A(N10634), .B(N10810));
NOR2XL inst_cellmath__198_0_I2797 (.Y(N10625), .A(N10810), .B(N44730));
NOR2XL inst_cellmath__198_0_I2798 (.Y(N10894), .A(N11027), .B(N10810));
NOR2XL inst_cellmath__198_0_I2799 (.Y(N10547), .A(N10810), .B(N10590));
NOR2XL inst_cellmath__198_0_I2800 (.Y(N10814), .A(N3809), .B(N10810));
NOR2XL inst_cellmath__198_0_I2801 (.Y(N10461), .A(N10973), .B(N10810));
NOR2XL inst_cellmath__198_0_I2802 (.Y(N10731), .A(N10810), .B(N10542));
NOR2XL inst_cellmath__198_0_I2803 (.Y(N11016), .A(N10810), .B(N10727));
NOR2XL inst_cellmath__198_0_I2804 (.Y(N10660), .A(N10810), .B(N10922));
NOR2XL inst_cellmath__198_0_I2805 (.Y(N10926), .A(N10491), .B(N10810));
OR2XL inst_cellmath__198_0_I2806 (.Y(N10452), .A(N10551), .B(N10810));
INVXL inst_cellmath__198_0_I2807 (.Y(N10962), .A(N10867));
NOR2XL inst_cellmath__198_0_I2808 (.Y(N10882), .A(N10431), .B(N10867));
NOR2XL inst_cellmath__198_0_I2809 (.Y(N10533), .A(N10634), .B(N10867));
NOR2XL inst_cellmath__198_0_I2810 (.Y(N10797), .A(N10867), .B(N44730));
NOR2XL inst_cellmath__198_0_I2811 (.Y(N10444), .A(N11027), .B(N10867));
NOR2XL inst_cellmath__198_0_I2812 (.Y(N10718), .A(N10867), .B(N10590));
NOR2XL inst_cellmath__198_0_I2813 (.Y(N11001), .A(N10867), .B(N3809));
NOR2XL inst_cellmath__198_0_I2814 (.Y(N10645), .A(N10973), .B(N10867));
NOR2XL inst_cellmath__198_0_I2815 (.Y(N10913), .A(N10867), .B(N10542));
NOR2XL inst_cellmath__198_0_I2816 (.Y(N10569), .A(N10867), .B(N10727));
NOR2XL inst_cellmath__198_0_I2817 (.Y(N10833), .A(N10867), .B(N10922));
NOR2XL inst_cellmath__198_0_I2818 (.Y(N10483), .A(N10491), .B(N10867));
OR2XL inst_cellmath__198_0_I2819 (.Y(N10598), .A(N10867), .B(N10551));
INVXL inst_cellmath__198_0_I2820 (.Y(N10517), .A(N10431));
NOR2XL inst_cellmath__198_0_I2821 (.Y(N10430), .A(N10431), .B(N10634));
NOR2XL inst_cellmath__198_0_I2822 (.Y(N10708), .A(N10431), .B(N44730));
NOR2XL inst_cellmath__198_0_I2823 (.Y(N10990), .A(N10431), .B(N11027));
NOR2XL inst_cellmath__198_0_I2824 (.Y(N10633), .A(N10431), .B(N10590));
NOR2X2 inst_cellmath__198_0_I2825 (.Y(N10902), .A(N3809), .B(N10431));
NOR2X1 inst_cellmath__198_0_I2826 (.Y(N10556), .A(N10973), .B(N10431));
NOR2X1 inst_cellmath__198_0_I2827 (.Y(N10822), .A(N10431), .B(N10542));
NOR2XL inst_cellmath__198_0_I2828 (.Y(N10469), .A(N10431), .B(N10727));
NOR2XL inst_cellmath__198_0_I2829 (.Y(N10739), .A(N10431), .B(N10922));
NOR2XL inst_cellmath__198_0_I2830 (.Y(N11026), .A(N10431), .B(N10491));
OR2XL inst_cellmath__198_0_I2831 (.Y(N10724), .A(N10431), .B(N10551));
INVXL inst_cellmath__198_0_I2832 (.Y(N10416), .A(N10634));
NOR2XL inst_cellmath__198_0_I2833 (.Y(N10972), .A(N10634), .B(N10823));
NOR2XL inst_cellmath__198_0_I2834 (.Y(N10620), .A(N10634), .B(N11027));
NOR2X1 inst_cellmath__198_0_I2835 (.Y(N10890), .A(N10634), .B(N10590));
NOR2X4 inst_cellmath__198_0_I2836 (.Y(N10541), .A(N10634), .B(N3809));
NOR2X4 inst_cellmath__198_0_I2837 (.Y(N10807), .A(N10634), .B(N10973));
NOR2XL inst_cellmath__198_0_I2838 (.Y(N10454), .A(N10634), .B(N10542));
NOR2XL inst_cellmath__198_0_I2839 (.Y(N10726), .A(N10634), .B(N10727));
NOR2XL inst_cellmath__198_0_I2840 (.Y(N11010), .A(N10634), .B(N10922));
NOR2XL inst_cellmath__198_0_I2841 (.Y(N10655), .A(N10634), .B(N10491));
OR2XL inst_cellmath__198_0_I2842 (.Y(N10862), .A(N10634), .B(N10551));
INVXL inst_cellmath__198_0_I2843 (.Y(N10683), .A(N44730));
NOR2X1 inst_cellmath__198_0_I2844 (.Y(N10609), .A(N10823), .B(N11027));
NOR2X2 inst_cellmath__198_0_I2845 (.Y(N10877), .A(N10590), .B(N10823));
NOR2X2 inst_cellmath__198_0_I2846 (.Y(N10528), .A(N3809), .B(N10823));
NOR2XL inst_cellmath__198_0_I2847 (.Y(N10792), .A(N10973), .B(N10823));
NOR2XL inst_cellmath__198_0_I2848 (.Y(N10439), .A(N10542), .B(N10823));
NOR2XL inst_cellmath__198_0_I2849 (.Y(N10715), .A(N10727), .B(N10823));
NOR2XL inst_cellmath__198_0_I2850 (.Y(N10996), .A(N10922), .B(N44730));
NOR2XL inst_cellmath__198_0_I2851 (.Y(N10640), .A(N10491), .B(N44730));
OR2XL inst_cellmath__198_0_I2852 (.Y(N11008), .A(N10551), .B(N44730));
INVX1 inst_cellmath__198_0_I2853 (.Y(N10671), .A(N11027));
NOR2X1 inst_cellmath__198_0_I2854 (.Y(N10597), .A(N10590), .B(N11027));
NOR2XL inst_cellmath__198_0_I2855 (.Y(N10860), .A(N11027), .B(N3809));
NOR2XL inst_cellmath__198_0_I2856 (.Y(N10512), .A(N11027), .B(N10973));
NOR2XL inst_cellmath__198_0_I2857 (.Y(N10776), .A(N11027), .B(N10542));
NOR2XL inst_cellmath__198_0_I2858 (.Y(N10424), .A(N11027), .B(N10727));
NOR2XL inst_cellmath__198_0_I2859 (.Y(N10702), .A(N11027), .B(N10922));
NOR2XL inst_cellmath__198_0_I2860 (.Y(N10981), .A(N11027), .B(N10491));
OR2XL inst_cellmath__198_0_I2861 (.Y(N10513), .A(N10551), .B(N11027));
INVX2 inst_cellmath__198_0_I2862 (.Y(N11019), .A(N10590));
NOR2XL inst_cellmath__198_0_I2863 (.Y(N10928), .A(N3809), .B(N10590));
NOR2XL inst_cellmath__198_0_I2864 (.Y(N10583), .A(N10973), .B(N10590));
NOR2XL inst_cellmath__198_0_I2865 (.Y(N10848), .A(N10542), .B(N10590));
NOR2XL inst_cellmath__198_0_I2866 (.Y(N10497), .A(N10727), .B(N10590));
NOR2XL inst_cellmath__198_0_I2867 (.Y(N10763), .A(N10922), .B(N10590));
NOR2XL inst_cellmath__198_0_I2868 (.Y(N10410), .A(N10491), .B(N10590));
OR2XL inst_cellmath__198_0_I2869 (.Y(N10653), .A(N10551), .B(N10590));
NOR2XL inst_cellmath__198_0_I2871 (.Y(N11005), .A(N3809), .B(N10973));
NOR2XL inst_cellmath__198_0_I2872 (.Y(N10649), .A(N3809), .B(N10542));
NOR2XL inst_cellmath__198_0_I2873 (.Y(N10917), .A(N3809), .B(N10727));
NOR2XL inst_cellmath__198_0_I2874 (.Y(N10573), .A(N3809), .B(N10922));
NOR2XL inst_cellmath__198_0_I2875 (.Y(N10838), .A(N3809), .B(N10491));
OR2XL inst_cellmath__198_0_I2876 (.Y(N10778), .A(N3809), .B(N10551));
INVXL inst_cellmath__198_0_I2877 (.Y(N10870), .A(N10973));
NOR2XL inst_cellmath__198_0_I2878 (.Y(N10786), .A(N10973), .B(N10542));
NOR2XL inst_cellmath__198_0_I2879 (.Y(N10433), .A(N10973), .B(N10727));
NOR2XL inst_cellmath__198_0_I2880 (.Y(N10710), .A(N10973), .B(N10922));
NOR2XL inst_cellmath__198_0_I2881 (.Y(N10992), .A(N10973), .B(N10491));
OR2XL inst_cellmath__198_0_I2882 (.Y(N10920), .A(N10551), .B(N10973));
INVXL inst_cellmath__198_0_I2883 (.Y(N11029), .A(N10542));
NOR2XL inst_cellmath__198_0_I2884 (.Y(N10936), .A(N10542), .B(N10727));
NOR2XL inst_cellmath__198_0_I2885 (.Y(N10592), .A(N10922), .B(N10542));
NOR2XL inst_cellmath__198_0_I2886 (.Y(N10855), .A(N10491), .B(N10542));
OR2XL inst_cellmath__198_0_I2887 (.Y(N10425), .A(N10551), .B(N10542));
INVXL inst_cellmath__198_0_I2888 (.Y(N10892), .A(N10727));
NOR2XL inst_cellmath__198_0_I2889 (.Y(N10809), .A(N10727), .B(N10922));
NOR2XL inst_cellmath__198_0_I2890 (.Y(N10457), .A(N10491), .B(N10727));
OR2XL inst_cellmath__198_0_I2891 (.Y(N10576), .A(N10551), .B(N10727));
INVXL inst_cellmath__198_0_I2892 (.Y(N10493), .A(N10922));
NOR2XL inst_cellmath__198_0_I2893 (.Y(N10403), .A(N10922), .B(N10491));
OR2XL inst_cellmath__198_0_I2894 (.Y(N10703), .A(N10922), .B(N10551));
INVXL inst_cellmath__198_0_I2895 (.Y(N10442), .A(N10491));
ADDHXL inst_cellmath__198_0_I2896 (.CO(N10984), .S(N10840), .A(N10481), .B(N10587));
INVXL inst_cellmath__198_0_I2897 (.Y(N11021), .A(N10840));
ADDHX1 inst_cellmath__198_0_I2898 (.CO(N10627), .S(N10489), .A(N10749), .B(N10852));
ADDHX1 inst_cellmath__198_0_I2899 (.CO(N10898), .S(N10756), .A(N10504), .B(N11037));
ADDFXL inst_cellmath__198_0_I2900 (.CO(N10550), .S(N10399), .A(N10953), .B(N10510), .CI(N10627));
ADDHX1 inst_cellmath__198_0_I2901 (.CO(N10817), .S(N10681), .A(N10676), .B(N10765));
ADDFX1 inst_cellmath__198_0_I2902 (.CO(N10465), .S(N10955), .A(N10898), .B(N10605), .CI(N10681));
ADDHX1 inst_cellmath__198_0_I2903 (.CO(N10734), .S(N10606), .A(N10947), .B(N10415));
ADDFX1 inst_cellmath__198_0_I2904 (.CO(N11020), .S(N10876), .A(N10962), .B(N10422), .CI(N10817));
ADDFXL inst_cellmath__198_0_I2905 (.CO(N10663), .S(N10525), .A(N10606), .B(N10874), .CI(N10465));
ADDHX1 inst_cellmath__198_0_I2906 (.CO(N10930), .S(N10789), .A(N10693), .B(N10600));
ADDFXL inst_cellmath__198_0_I2907 (.CO(N10585), .S(N10438), .A(N10523), .B(N10699), .CI(N10734));
ADDFXL inst_cellmath__198_0_I2908 (.CO(N10850), .S(N10714), .A(N11020), .B(N10789), .CI(N10438));
ADDHX1 inst_cellmath__198_0_I2909 (.CO(N10500), .S(N10995), .A(N10865), .B(N10970));
ADDFXL inst_cellmath__198_0_I2910 (.CO(N10764), .S(N10639), .A(N10517), .B(N10979), .CI(N10882));
ADDFX1 inst_cellmath__198_0_I2911 (.CO(N10412), .S(N10909), .A(N10995), .B(N10788), .CI(N10930));
ADDFXL inst_cellmath__198_0_I2912 (.CO(N10691), .S(N10561), .A(N10639), .B(N10585), .CI(N10909));
ADDHX1 inst_cellmath__198_0_I2913 (.CO(N10967), .S(N10829), .A(N10516), .B(N10619));
ADDFX1 inst_cellmath__198_0_I2914 (.CO(N10617), .S(N10477), .A(N10533), .B(N10625), .CI(N10500));
ADDFXL inst_cellmath__198_0_I2915 (.CO(N10885), .S(N10743), .A(N10436), .B(N10829), .CI(N10764));
ADDFXL inst_cellmath__198_0_I2916 (.CO(N10536), .S(N11033), .A(N10412), .B(N10477), .CI(N10743));
ADDHX1 inst_cellmath__198_0_I2917 (.CO(N10801), .S(N10670), .A(N10781), .B(N10416));
ADDFX1 inst_cellmath__198_0_I2918 (.CO(N10449), .S(N10940), .A(N10889), .B(N10430), .CI(N10894));
ADDFX1 inst_cellmath__198_0_I2919 (.CO(N10720), .S(N10596), .A(N10967), .B(N10797), .CI(N10670));
ADDFX1 inst_cellmath__198_0_I2920 (.CO(N11006), .S(N10858), .A(N10712), .B(N10617), .CI(N10940));
ADDFXL inst_cellmath__198_0_I2921 (.CO(N10651), .S(N10511), .A(N10596), .B(N10885), .CI(N10858));
ADDHXL inst_cellmath__198_0_I2922 (.CO(N10918), .S(N10775), .A(N10428), .B(N10538));
ADDFXL inst_cellmath__198_0_I2923 (.CO(N10574), .S(N10423), .A(N10547), .B(N10708), .CI(N10801));
ADDFX1 inst_cellmath__198_0_I2924 (.CO(N10839), .S(N10700), .A(N10994), .B(N10444), .CI(N10775));
ADDFX1 inst_cellmath__198_0_I2925 (.CO(N10487), .S(N10980), .A(N10720), .B(N10449), .CI(N10423));
ADDFX1 inst_cellmath__198_0_I2926 (.CO(N10753), .S(N10626), .A(N11006), .B(N10700), .CI(N10980));
ADDHXL inst_cellmath__198_0_I2927 (.CO(N10398), .S(N10895), .A(N10972), .B(N10706));
ADDFX1 inst_cellmath__198_0_I2928 (.CO(N10679), .S(N10548), .A(N10990), .B(N10683), .CI(N10804));
ADDFXL inst_cellmath__198_0_I2929 (.CO(N10951), .S(N10815), .A(N10718), .B(N10814), .CI(N10918));
ADDFXL inst_cellmath__198_0_I2930 (.CO(N10604), .S(N10462), .A(N10895), .B(N10637), .CI(N10574));
ADDFX1 inst_cellmath__198_0_I2931 (.CO(N10872), .S(N10732), .A(N10839), .B(N10548), .CI(N10815));
ADDFX1 inst_cellmath__198_0_I2932 (.CO(N10520), .S(N11017), .A(N10487), .B(N10462), .CI(N10732));
ADDHX1 inst_cellmath__198_0_I2933 (.CO(N10787), .S(N10661), .A(N10987), .B(N10620));
ADDFX1 inst_cellmath__198_0_I2934 (.CO(N10434), .S(N10927), .A(N10451), .B(N10633), .CI(N10461));
ADDFXL inst_cellmath__198_0_I2935 (.CO(N10711), .S(N10582), .A(N11001), .B(N10907), .CI(N10398));
ADDFXL inst_cellmath__198_0_I2937 (.CO(N10636), .S(N10496), .A(N10582), .B(N10927), .CI(N10604));
ADDFX1 inst_cellmath__198_0_I29683 (.CO(N45620), .S(N10847), .A(N10679), .B(N10661), .CI(N10951));
ADDFXL inst_cellmath__198_0_I2938 (.CO(N10906), .S(N10761), .A(N10847), .B(N10872), .CI(N10496));
ADDHXL inst_cellmath__198_0_I2939 (.CO(N10558), .S(N10408), .A(N10890), .B(N10609));
ADDFXL inst_cellmath__198_0_I2940 (.CO(N10825), .S(N10688), .A(N10630), .B(N10671), .CI(N10902));
ADDFXL inst_cellmath__198_0_I29686 (.CO(N45575), .S(N10883), .A(N10434), .B(N10688), .CI(N10711));
ADDFXL inst_cellmath__198_0_I29685 (.CO(N45611), .S(N45598), .A(N10787), .B(N10560), .CI(N10408));
ADDFX1 inst_cellmath__198_0_I29684 (.CO(N45583), .S(N45569), .A(N10731), .B(N10722), .CI(N10645));
ADDFX1 inst_cellmath__198_0_I29687 (.CO(N45604), .S(N10534), .A(N45598), .B(N45569), .CI(N45620));
ADDFHX1 inst_cellmath__198_0_I2945 (.CO(N10937), .S(N10798), .A(N10636), .B(N10883), .CI(N10534));
INVX1 xnor2_A_I30579 (.Y(N45774), .A(N10541));
MXI2XL xnor2_A_I30580 (.Y(N10445), .A(N10541), .B(N45774), .S0(N10877));
OR2XL inst_cellmath__198_0_I2947 (.Y(N10593), .A(N10877), .B(N10541));
ADDFHXL inst_cellmath__198_0_I2954 (.CO(N10893), .S(N10750), .A(N11019), .B(N10807), .CI(N10528));
ADDFXL inst_cellmath__198_0_I2961 (.CO(N10925), .S(N10784), .A(N10454), .B(N10469), .CI(N10792));
ADDFX1 inst_cellmath__198_0_I2962 (.CO(N10581), .S(N10432), .A(N10860), .B(N10926), .CI(N10833));
ADDFXL inst_cellmath__198_0_I29694 (.CO(N10544), .S(N45592), .A(N10822), .B(N10597), .CI(N10805));
ADDFHXL inst_cellmath__198_0_I2963 (.CO(N10845), .S(N10709), .A(N10893), .B(N10944), .CI(N10544));
ADDFX1 inst_cellmath__198_0_I29695 (.CO(N10811), .S(N45621), .A(N10660), .B(N10593), .CI(N10569));
ADDFX1 inst_cellmath__198_0_I2964 (.CO(N10495), .S(N10991), .A(N10811), .B(N10784), .CI(N10432));
ADDFX1 inst_cellmath__198_0_I29688 (.CO(N45631), .S(N45618), .A(N11007), .B(N10556), .CI(N10673));
ADDFHXL inst_cellmath__198_0_I29696 (.CO(N10458), .S(N45584), .A(N45631), .B(N10476), .CI(N10750));
ADDFHX1 inst_cellmath__198_0_I29689 (.CO(N45595), .S(N45581), .A(N11016), .B(N10913), .CI(N10558));
ADDFXL inst_cellmath__198_0_I29690 (.CO(N45624), .S(N45608), .A(N10827), .B(N10445), .CI(N10825));
ADDFHXL inst_cellmath__198_0_I29697 (.CO(N10729), .S(N45612), .A(N45595), .B(N45592), .CI(N45624));
ADDFHXL inst_cellmath__198_0_I2965 (.CO(N10759), .S(N10635), .A(N10709), .B(N10458), .CI(N10729));
ADDFX1 inst_cellmath__198_0_I29691 (.CO(N45587), .S(N45572), .A(N45618), .B(N45583), .CI(N45611));
ADDFHXL inst_cellmath__198_0_I29698 (.CO(N11013), .S(N45576), .A(N45584), .B(N45621), .CI(N45587));
ADDFHXL inst_cellmath__198_0_I2966 (.CO(N10406), .S(N10903), .A(N11013), .B(N10991), .CI(N10635));
ADDFXL inst_cellmath__198_0_I2967 (.CO(N10686), .S(N10557), .A(N3810), .B(N10928), .CI(N10439));
ADDFXL inst_cellmath__198_0_I2968 (.CO(N10960), .S(N10824), .A(N10726), .B(N10512), .CI(N10739));
ADDFXL inst_cellmath__198_0_I2969 (.CO(N10613), .S(N10470), .A(N10483), .B(N10452), .CI(N10925));
ADDFX1 inst_cellmath__198_0_I2970 (.CO(N10881), .S(N10740), .A(N10581), .B(N10557), .CI(N10824));
ADDFXL inst_cellmath__198_0_I2971 (.CO(N10530), .S(N11028), .A(N10470), .B(N10845), .CI(N10495));
ADDFHXL inst_cellmath__198_0_I2972 (.CO(N10796), .S(N10667), .A(N10740), .B(N10759), .CI(N11028));
ADDFX1 inst_cellmath__198_0_I2973 (.CO(N10443), .S(N10935), .A(N10583), .B(N11026), .CI(N10715));
ADDFX1 inst_cellmath__198_0_I2974 (.CO(N10717), .S(N10591), .A(N11010), .B(N10776), .CI(N10598));
ADDFX1 inst_cellmath__198_0_I2975 (.CO(N11000), .S(N10853), .A(N10960), .B(N10686), .CI(N10935));
ADDFHXL inst_cellmath__198_0_I2976 (.CO(N10644), .S(N10505), .A(N10613), .B(N10591), .CI(N10881));
ADDFHX1 inst_cellmath__198_0_I2977 (.CO(N10911), .S(N10768), .A(N10853), .B(N10530), .CI(N10505));
ADDFXL inst_cellmath__198_0_I2978 (.CO(N10566), .S(N10417), .A(N10870), .B(N10655), .CI(N11005));
ADDFX1 inst_cellmath__198_0_I2979 (.CO(N10832), .S(N10694), .A(N10424), .B(N10848), .CI(N10724));
ADDFX1 inst_cellmath__198_0_I2980 (.CO(N10480), .S(N10974), .A(N10996), .B(N10443), .CI(N10417));
ADDFHXL inst_cellmath__198_0_I2981 (.CO(N10748), .S(N10621), .A(N10694), .B(N10717), .CI(N11000));
ADDFXL inst_cellmath__198_0_I2982 (.CO(N11038), .S(N10891), .A(N10644), .B(N10974), .CI(N10621));
ADDFX1 inst_cellmath__198_0_I2983 (.CO(N10675), .S(N10543), .A(N10649), .B(N10640), .CI(N10497));
ADDFXL inst_cellmath__198_0_I2984 (.CO(N10946), .S(N10808), .A(N10702), .B(N10862), .CI(N10566));
ADDFXL inst_cellmath__198_0_I2985 (.CO(N10601), .S(N10455), .A(N10543), .B(N10832), .CI(N10480));
ADDFXL inst_cellmath__198_0_I2986 (.CO(N10864), .S(N10728), .A(N10748), .B(N10808), .CI(N10455));
ADDFX1 inst_cellmath__198_0_I2987 (.CO(N10515), .S(N11011), .A(N11029), .B(N10786), .CI(N10917));
ADDFX1 inst_cellmath__198_0_I2988 (.CO(N10782), .S(N10656), .A(N10981), .B(N10763), .CI(N11008));
ADDFX1 inst_cellmath__198_0_I2989 (.CO(N10427), .S(N10923), .A(N11011), .B(N10675), .CI(N10946));
ADDFXL inst_cellmath__198_0_I2990 (.CO(N10705), .S(N10579), .A(N10601), .B(N10656), .CI(N10923));
ADDFX1 inst_cellmath__198_0_I2991 (.CO(N10988), .S(N10842), .A(N10433), .B(N10410), .CI(N10573));
ADDFX1 inst_cellmath__198_0_I2992 (.CO(N10629), .S(N10492), .A(N10515), .B(N10513), .CI(N10782));
ADDFX1 inst_cellmath__198_0_I2993 (.CO(N10900), .S(N10758), .A(N10427), .B(N10842), .CI(N10492));
ADDFX1 inst_cellmath__198_0_I2994 (.CO(N10554), .S(N10401), .A(N10838), .B(N10892), .CI(N10936));
ADDFX1 inst_cellmath__198_0_I2995 (.CO(N10819), .S(N10684), .A(N10710), .B(N10653), .CI(N10988));
ADDFX1 inst_cellmath__198_0_I2996 (.CO(N10468), .S(N10958), .A(N10629), .B(N10401), .CI(N10684));
ADDFX1 inst_cellmath__198_0_I2997 (.CO(N10737), .S(N10610), .A(N10778), .B(N10992), .CI(N10592));
ADDFX1 inst_cellmath__198_0_I2998 (.CO(N11023), .S(N10880), .A(N10610), .B(N10554), .CI(N10819));
ADDFX1 inst_cellmath__198_0_I2999 (.CO(N10666), .S(N10529), .A(N10493), .B(N10855), .CI(N10920));
ADDFX1 inst_cellmath__198_0_I3000 (.CO(N10933), .S(N10793), .A(N10737), .B(N10809), .CI(N10529));
ADDFX1 inst_cellmath__198_0_I3001 (.CO(N10586), .S(N10441), .A(N10425), .B(N10457), .CI(N10666));
ADDFX1 inst_cellmath__198_0_I3002 (.CO(N10851), .S(N10716), .A(N10403), .B(N10442), .CI(N10576));
NAND2XL inst_cellmath__198_0_I3005 (.Y(N10414), .A(N10984), .B(N10489));
AND2XL inst_cellmath__198_0_I3007 (.Y(N10692), .A(N10756), .B(N10399));
NAND2XL inst_cellmath__198_0_I3009 (.Y(N10969), .A(N10550), .B(N10955));
OR2XL inst_cellmath__198_0_I3010 (.Y(N10479), .A(N10876), .B(N10525));
AND2XL inst_cellmath__198_0_I3011 (.Y(N10618), .A(N10876), .B(N10525));
NOR2XL inst_cellmath__198_0_I3012 (.Y(N10745), .A(N10663), .B(N10714));
NAND2X1 inst_cellmath__198_0_I3013 (.Y(N10888), .A(N10663), .B(N10714));
NOR2X1 inst_cellmath__198_0_I3014 (.Y(N11035), .A(N10850), .B(N10561));
NOR2XL inst_cellmath__198_0_I3016 (.Y(N10672), .A(N10691), .B(N11033));
NAND2X2 inst_cellmath__198_0_I3017 (.Y(N10803), .A(N10691), .B(N11033));
NOR2XL inst_cellmath__198_0_I3018 (.Y(N10942), .A(N10536), .B(N10511));
NAND2X1 inst_cellmath__198_0_I3019 (.Y(N10450), .A(N10536), .B(N10511));
NOR3XL inst_cellmath__198_0_I11212 (.Y(N10861), .A(N10418), .B(N10622), .C(N10878));
NOR2XL inst_cellmath__198_0_I3023 (.Y(N10790), .A(N10622), .B(N11021));
OAI2BB2XL inst_cellmath__198_0_I10715 (.Y(N10982), .A0N(N10622), .A1N(N11021), .B0(N10861), .B1(N10790));
AOI2BB2X1 inst_cellmath__198_0_I10716 (.Y(N10816), .A0N(N10984), .A1N(N10489), .B0(N10982), .B1(N10414));
OAI22X1 inst_cellmath__198_0_I10717 (.Y(N10584), .A0(N10692), .A1(N10816), .B0(N10756), .B1(N10399));
AOI2BB2X1 inst_cellmath__198_0_I10718 (.Y(N10966), .A0N(N10550), .A1N(N10955), .B0(N10584), .B1(N10969));
OAI21X1 inst_cellmath__198_0_I3033 (.Y(N10650), .A0(N10618), .A1(N10966), .B0(N10479));
AOI21X2 inst_cellmath__198_0_I3034 (.Y(N10950), .A0(N10888), .A1(N10650), .B0(N10745));
AOI21X2 inst_cellmath__198_0_I3035 (.Y(N10871), .A0(N11035), .A1(N10803), .B0(N10672));
OAI2BB1X1 inst_cellmath__198_0_I10722 (.Y(N11015), .A0N(N10850), .A1N(N10561), .B0(N10803));
OAI21X2 inst_cellmath__198_0_I3037 (.Y(N10472), .A0(N11015), .A1(N10950), .B0(N10871));
AOI21X2 inst_cellmath__198_0_I3040 (.Y(N10975), .A0(N10450), .A1(N10472), .B0(N10942));
INVX1 inst_cellmath__198_0_I3061 (.Y(N10747), .A(N10975));
NOR2XL inst_cellmath__198_0_I3062 (.Y(N11036), .A(N10651), .B(N10626));
NAND2X1 inst_cellmath__198_0_I3063 (.Y(N10540), .A(N10651), .B(N10626));
NOR2X1 inst_cellmath__198_0_I3064 (.Y(N10674), .A(N10753), .B(N11017));
NOR2XL inst_cellmath__198_0_I3066 (.Y(N10945), .A(N10520), .B(N10761));
NAND2X2 inst_cellmath__198_0_I3067 (.Y(N10453), .A(N10520), .B(N10761));
NOR2X2 inst_cellmath__198_0_I3068 (.Y(N10599), .A(N10906), .B(N10798));
NAND2X2 inst_cellmath__198_0_I3069 (.Y(N10725), .A(N10906), .B(N10798));
ADDFXL inst_cellmath__198_0_I29692 (.CO(N45615), .S(N45601), .A(N45581), .B(N45608), .CI(N45575));
ADDFHX1 inst_cellmath__198_0_I29693 (.CO(N10623), .S(N10484), .A(N45604), .B(N45572), .CI(N45601));
NOR2X1 inst_cellmath__198_0_I3070 (.Y(N10863), .A(N10937), .B(N10484));
NAND2X4 inst_cellmath__198_0_I3071 (.Y(N11009), .A(N10937), .B(N10484));
ADDFHXL inst_cellmath__198_0_I29699 (.CO(N10658), .S(N10518), .A(N45615), .B(N45612), .CI(N45576));
NOR2X2 inst_cellmath__198_0_I3072 (.Y(N10514), .A(N10623), .B(N10518));
NAND2X2 inst_cellmath__198_0_I29700 (.Y(N10654), .A(N10623), .B(N10518));
NOR2X1 inst_cellmath__198_0_I3074 (.Y(N10780), .A(N10658), .B(N10903));
NAND2X4 inst_cellmath__198_0_I3075 (.Y(N10921), .A(N10658), .B(N10903));
NOR2X2 inst_cellmath__198_0_I3076 (.Y(N10426), .A(N10406), .B(N10667));
NAND2X2 inst_cellmath__198_0_I3077 (.Y(N10577), .A(N10406), .B(N10667));
NOR2X1 inst_cellmath__198_0_I3078 (.Y(N10704), .A(N10796), .B(N10768));
NAND2X4 inst_cellmath__198_0_I3079 (.Y(N10841), .A(N10796), .B(N10768));
NOR2X1 inst_cellmath__198_0_I3080 (.Y(N10986), .A(N10911), .B(N10891));
NAND2X2 inst_cellmath__198_0_I3081 (.Y(N10490), .A(N10911), .B(N10891));
NOR2XL inst_cellmath__198_0_I3082 (.Y(N10628), .A(N11038), .B(N10728));
NAND2X2 inst_cellmath__198_0_I3083 (.Y(N10757), .A(N11038), .B(N10728));
NOR2XL inst_cellmath__198_0_I3086 (.Y(N10552), .A(N10758), .B(N10705));
NAND2X1 inst_cellmath__198_0_I3087 (.Y(N10682), .A(N10758), .B(N10705));
NOR2XL inst_cellmath__198_0_I3088 (.Y(N10818), .A(N10900), .B(N10958));
NAND2XL inst_cellmath__198_0_I3089 (.Y(N10957), .A(N10900), .B(N10958));
NOR2XL inst_cellmath__198_0_I3090 (.Y(N10467), .A(N10468), .B(N10880));
NAND2XL inst_cellmath__198_0_I3091 (.Y(N10608), .A(N10468), .B(N10880));
NOR2XL inst_cellmath__198_0_I3092 (.Y(N10736), .A(N10793), .B(N11023));
NAND2XL inst_cellmath__198_0_I3093 (.Y(N10879), .A(N10793), .B(N11023));
NOR2XL inst_cellmath__198_0_I3094 (.Y(N11022), .A(N10933), .B(N10441));
NAND2XL inst_cellmath__198_0_I3095 (.Y(N10527), .A(N10933), .B(N10441));
NOR2XL inst_cellmath__198_0_I3096 (.Y(N10665), .A(N10716), .B(N10586));
NAND2XL inst_cellmath__198_0_I3097 (.Y(N10791), .A(N10716), .B(N10586));
NOR2XL inst_cellmath__198_0_I3098 (.Y(N10932), .A(N10703), .B(N10851));
NAND2XL inst_cellmath__198_0_I3099 (.Y(N10440), .A(N10703), .B(N10851));
AOI21X2 inst_cellmath__198_0_I3100 (.Y(N10502), .A0(N10540), .A1(N10747), .B0(N11036));
AOI21X2 inst_cellmath__198_0_I3101 (.Y(N10413), .A0(N10453), .A1(N10674), .B0(N10945));
OAI2BB1X1 inst_cellmath__198_0_I10727 (.Y(N10562), .A0N(N10753), .A1N(N11017), .B0(N10453));
AOI21X4 inst_cellmath__198_0_I3103 (.Y(N10968), .A0(N11009), .A1(N10599), .B0(N10863));
NAND2X2 inst_cellmath__198_0_I3104 (.Y(N10478), .A(N11009), .B(N10725));
AOI21X4 inst_cellmath__198_0_I3105 (.Y(N10887), .A0(N10921), .A1(N10514), .B0(N10780));
NAND2X2 inst_cellmath__198_0_I3106 (.Y(N11034), .A(N10921), .B(N10654));
AOI21X4 inst_cellmath__198_0_I3107 (.Y(N10802), .A0(N10426), .A1(N10841), .B0(N10704));
NAND2X4 inst_cellmath__198_0_I3108 (.Y(N10941), .A(N10841), .B(N10577));
AOI21X2 inst_cellmath__198_0_I3109 (.Y(N10721), .A0(N10757), .A1(N10986), .B0(N10628));
NAND2X4 inst_cellmath__198_0_I3110 (.Y(N10859), .A(N10757), .B(N10490));
NOR2X1 inst_cellmath__203_0_I29529 (.Y(N10899), .A(N10864), .B(N10579));
AOI21X1 inst_cellmath__198_0_I3111 (.Y(N10652), .A0(N10682), .A1(N10899), .B0(N10552));
NAND2X1 inst_cellmath__203_0_I29530 (.Y(N10400), .A(N10864), .B(N10579));
NAND2XL inst_cellmath__198_0_I3112 (.Y(N10777), .A(N10682), .B(N10400));
INVXL inst_cellmath__198_0_I3113 (.Y(N10475), .A(N10818));
INVXL inst_cellmath__198_0_I3114 (.Y(N10616), .A(N10957));
AOI21XL inst_cellmath__198_0_I3115 (.Y(N10575), .A0(N10608), .A1(N10818), .B0(N10467));
NAND2XL inst_cellmath__198_0_I3116 (.Y(N10701), .A(N10608), .B(N10957));
OAI21XL inst_cellmath__198_0_I3117 (.Y(N10754), .A0(N10616), .A1(N10652), .B0(N10475));
AOI21XL inst_cellmath__198_0_I3118 (.Y(N10952), .A0(N10527), .A1(N10736), .B0(N11022));
NAND2XL inst_cellmath__198_0_I3119 (.Y(N10463), .A(N10527), .B(N10879));
INVXL inst_cellmath__198_0_I3120 (.Y(N10939), .A(N10665));
INVXL inst_cellmath__198_0_I3121 (.Y(N10447), .A(N10791));
AOI21XL inst_cellmath__198_0_I3122 (.Y(N10873), .A0(N10440), .A1(N10665), .B0(N10932));
NAND2XL inst_cellmath__198_0_I3123 (.Y(N11018), .A(N10440), .B(N10791));
OAI21XL inst_cellmath__198_0_I3124 (.Y(N10435), .A0(N10447), .A1(N10952), .B0(N10939));
OA21XL inst_cellmath__198_0_I3125 (.Y(N10698), .A0(N10701), .A1(N10652), .B0(N10575));
OR2XL inst_cellmath__198_0_I3126 (.Y(N10836), .A(N10701), .B(N10777));
OA21X1 inst_cellmath__198_0_I3127 (.Y(N10545), .A0(N11018), .A1(N10952), .B0(N10873));
OR2XL inst_cellmath__198_0_I3128 (.Y(N10678), .A(N11018), .B(N10463));
INVXL inst_cellmath__198_0_I3129 (.Y(N10812), .A(N10502));
OAI21X2 inst_cellmath__198_0_I3130 (.Y(N10595), .A0(N10562), .A1(N10502), .B0(N10413));
OAI21X2 inst_cellmath__198_0_I3131 (.Y(N10857), .A0(N10478), .A1(N10413), .B0(N10968));
NOR2X1 inst_cellmath__198_0_I3132 (.Y(N11004), .A(N10562), .B(N10478));
OAI21X2 inst_cellmath__198_0_I3133 (.Y(N10509), .A0(N10968), .A1(N11034), .B0(N10887));
NOR2X2 inst_cellmath__198_0_I3134 (.Y(N10648), .A(N10478), .B(N11034));
OAI21X2 inst_cellmath__198_0_I3135 (.Y(N10773), .A0(N10941), .A1(N10887), .B0(N10802));
NOR2X2 inst_cellmath__198_0_I3136 (.Y(N10916), .A(N10941), .B(N11034));
OAI21X2 inst_cellmath__198_0_I3137 (.Y(N10421), .A0(N10859), .A1(N10802), .B0(N10721));
NOR2X2 inst_cellmath__198_0_I3138 (.Y(N10572), .A(N10859), .B(N10941));
OAI21XL inst_cellmath__198_0_I3139 (.Y(N10697), .A0(N10836), .A1(N10721), .B0(N10698));
NOR2XL inst_cellmath__198_0_I3140 (.Y(N10837), .A(N10836), .B(N10859));
OAI21XL inst_cellmath__198_0_I3141 (.Y(N10978), .A0(N10678), .A1(N10698), .B0(N10545));
NOR2XL inst_cellmath__198_0_I3142 (.Y(N10486), .A(N10678), .B(N10836));
INVXL inst_cellmath__198_0_I3143 (.Y(N10949), .A(N10812));
AOI21X2 inst_cellmath__198_0_I3145 (.Y(N10546), .A0(N11004), .A1(N10812), .B0(N10857));
AOI21X1 inst_cellmath__198_0_I3146 (.Y(N10813), .A0(N10648), .A1(N10595), .B0(N10509));
AOI21X1 inst_cellmath__198_0_I3147 (.Y(N10459), .A0(N10916), .A1(N10857), .B0(N10773));
NAND2X1 inst_cellmath__198_0_I3148 (.Y(N10603), .A(N11004), .B(N10916));
AOI21X1 inst_cellmath__198_0_I3151 (.Y(N11014), .A0(N10837), .A1(N10773), .B0(N10697));
NAND2X1 inst_cellmath__198_0_I3152 (.Y(N10519), .A(N10837), .B(N10916));
AOI21XL inst_cellmath__198_0_I3153 (.Y(N10659), .A0(N10486), .A1(N10421), .B0(N10978));
NAND2XL inst_cellmath__198_0_I3154 (.Y(N10785), .A(N10486), .B(N10572));
OAI21X1 inst_cellmath__198_0_I3155 (.Y(N10760), .A0(N10949), .A1(N10603), .B0(N10459));
OAI21X2 inst_cellmath__198_0_I3157 (.Y(N10687), .A0(N10519), .A1(N10546), .B0(N11014));
OAI21XL inst_cellmath__198_0_I3158 (.Y(N10961), .A0(N10785), .A1(N10813), .B0(N10659));
INVXL inst_cellmath__198_0_I3160 (.Y(N10471), .A(N10952));
NAND2BXL inst_cellmath__198_0_I3165 (.Y(N10843), .AN(N10863), .B(N11009));
NAND2BXL inst_cellmath__198_0_I3166 (.Y(N10631), .AN(N10514), .B(N10654));
NAND2BXL inst_cellmath__198_0_I3167 (.Y(N10402), .AN(N10780), .B(N10921));
NAND2BXL inst_cellmath__198_0_I3168 (.Y(N10820), .AN(N10426), .B(N10577));
NAND2BXL inst_cellmath__198_0_I3169 (.Y(N10611), .AN(N10704), .B(N10841));
NAND2BXL inst_cellmath__198_0_I3170 (.Y(N11024), .AN(N10986), .B(N10490));
NAND2BXL inst_cellmath__198_0_I3171 (.Y(N10794), .AN(N10628), .B(N10757));
NAND2BXL inst_cellmath__198_0_I3172 (.Y(N10588), .AN(N10899), .B(N10400));
NAND2BXL inst_cellmath__198_0_I3175 (.Y(N10565), .AN(N10467), .B(N10608));
NAND2BXL inst_cellmath__198_0_I3176 (.Y(N10971), .AN(N10736), .B(N10879));
NAND2BXL inst_cellmath__198_0_I3177 (.Y(N10746), .AN(N11022), .B(N10527));
NAND2BXL inst_cellmath__198_0_I3178 (.Y(N10539), .AN(N10665), .B(N10791));
NAND2BXL inst_cellmath__198_0_I3179 (.Y(N10943), .AN(N10932), .B(N10440));
NAND2XL inst_cellmath__198_0_I3180 (.Y(N10723), .A(N10491), .B(inst_cellmath__115__W1[0]));
XNOR2X1 inst_cellmath__198_0_I3184 (.Y(inst_cellmath__198[18]), .A(N10631), .B(N10546));
XNOR2X1 inst_cellmath__198_0_I3185 (.Y(inst_cellmath__198[20]), .A(N10820), .B(N10813));
INVXL xnor2_A_I30581 (.Y(N45780), .A(N11024));
MXI2XL xnor2_A_I30582 (.Y(inst_cellmath__198[22]), .A(N11024), .B(N45780), .S0(N10760));
NAND2X2 inst_cellmath__203_0_I29533 (.Y(N45208), .A(N10572), .B(N10648));
INVX1 inst_cellmath__203_0_I29531 (.Y(N10460), .A(N10595));
AOI21X2 inst_cellmath__203_0_I29532 (.Y(N45200), .A0(N10572), .A1(N10509), .B0(N10421));
OAI21X4 inst_cellmath__203_0_I29665 (.Y(N10407), .A0(N45208), .A1(N10460), .B0(N45200));
XNOR2X1 inst_cellmath__198_0_I3187 (.Y(inst_cellmath__198[24]), .A(N10588), .B(N10407));
XNOR2X1 inst_cellmath__198_0_I3188 (.Y(inst_cellmath__198[28]), .A(N10971), .B(N10687));
XNOR2XL inst_cellmath__198_0_I3189 (.Y(inst_cellmath__198[32]), .A(N10723), .B(N10961));
INVXL xnor2_A_I30583 (.Y(N45786), .A(N10725));
MXI2XL xnor2_A_I30584 (.Y(N10755), .A(N10725), .B(N45786), .S0(N10843));
INVXL xnor2_A_I30585 (.Y(N45792), .A(N10599));
MXI2XL xnor2_A_I30586 (.Y(N10897), .A(N10599), .B(N45792), .S0(N10843));
XNOR2X1 inst_cellmath__198_0_I3196 (.Y(N10549), .A(N10654), .B(N10402));
XNOR2X1 inst_cellmath__198_0_I3197 (.Y(N10680), .A(N10514), .B(N10402));
MXI2X1 inst_cellmath__198_0_I3198 (.Y(inst_cellmath__198[19]), .A(N10549), .B(N10680), .S0(N10546));
XNOR2X1 inst_cellmath__198_0_I3199 (.Y(N10954), .A(N10577), .B(N10611));
XNOR2X1 inst_cellmath__198_0_I3200 (.Y(N10464), .A(N10426), .B(N10611));
MX2X1 inst_cellmath__198_0_I3201 (.Y(inst_cellmath__198[21]), .A(N10954), .B(N10464), .S0(N10813));
XNOR2X1 inst_cellmath__198_0_I3202 (.Y(N10733), .A(N10794), .B(N10490));
XNOR2X1 inst_cellmath__198_0_I3203 (.Y(N10875), .A(N10794), .B(N10986));
MX2XL inst_cellmath__198_0_I3204 (.Y(inst_cellmath__198[23]), .A(N10875), .B(N10733), .S0(N10760));
BUFX2 inst_cellmath__198_0_I10728 (.Y(N23282), .A(inst_cellmath__198[23]));
XNOR2X1 inst_cellmath__198_0_I3212 (.Y(N10713), .A(N10565), .B(N10754));
NOR2XL inst_cellmath__198_0_I3213 (.Y(N10854), .A(N10616), .B(N10777));
NOR2XL inst_cellmath__198_0_I3214 (.Y(N10498), .A(N10854), .B(N10754));
XOR2XL inst_cellmath__198_0_I3215 (.Y(N10849), .A(N10565), .B(N10498));
MX2XL inst_cellmath__198_0_I3216 (.Y(inst_cellmath__198[27]), .A(N10713), .B(N10849), .S0(N10407));
XNOR2X1 inst_cellmath__198_0_I3217 (.Y(N10499), .A(N10746), .B(N10879));
XNOR2X1 inst_cellmath__198_0_I3218 (.Y(N10638), .A(N10746), .B(N10736));
MX2XL inst_cellmath__198_0_I3219 (.Y(inst_cellmath__198[29]), .A(N10638), .B(N10499), .S0(N10687));
XNOR2X1 inst_cellmath__198_0_I3220 (.Y(N10908), .A(N10539), .B(N10471));
NOR2BX1 inst_cellmath__198_0_I3221 (.Y(N10800), .AN(N10463), .B(N10471));
XOR2XL inst_cellmath__198_0_I3222 (.Y(N10411), .A(N10539), .B(N10800));
MX2X1 inst_cellmath__198_0_I3223 (.Y(inst_cellmath__198[30]), .A(N10908), .B(N10411), .S0(N10687));
XNOR2X1 inst_cellmath__198_0_I3224 (.Y(N10690), .A(N10943), .B(N10435));
NOR2XL inst_cellmath__198_0_I3225 (.Y(N10568), .A(N10447), .B(N10463));
NOR2XL inst_cellmath__198_0_I3226 (.Y(N10774), .A(N10568), .B(N10435));
XOR2XL inst_cellmath__198_0_I3227 (.Y(N10828), .A(N10943), .B(N10774));
MXI2X1 inst_cellmath__198_0_I3228 (.Y(inst_cellmath__198[31]), .A(N10690), .B(N10828), .S0(N10687));
NAND3XL hyperpropagate_4_1_A_I11460 (.Y(N23367), .A(N8990), .B(N8933), .C(N8003));
NOR2XL hyperpropagate_4_1_A_I11461 (.Y(N12104), .A(N8540), .B(N23367));
INVXL inst_cellmath__203_0_I3230 (.Y(N12468), .A(inst_cellmath__197[1]));
NOR4X1 inst_cellmath__203_0_I10993 (.Y(N12807), .A(N8982), .B(N7948), .C(N8374), .D(N9032));
INVXL inst_cellmath__203_0_I3232 (.Y(N13175), .A(inst_cellmath__197[3]));
NAND3XL hyperpropagate_4_1_A_I11462 (.Y(N23375), .A(N8872), .B(N8594), .C(N8390));
NOR2XL hyperpropagate_4_1_A_I11463 (.Y(N11881), .A(N9122), .B(N23375));
INVX1 inst_cellmath__203_0_I3234 (.Y(N12253), .A(inst_cellmath__197[5]));
INVX1 inst_cellmath__203_0_I3235 (.Y(N12618), .A(inst_cellmath__197[6]));
NOR4X1 inst_cellmath__203_0_I11219 (.Y(N12956), .A(N8805), .B(N8733), .C(N8045), .D(N8376));
NOR4BX1 inst_cellmath__203_0_I11220 (.Y(N13340), .AN(N8838), .B(N8622), .C(N8707), .D(N8497));
NOR3BX1 inst_cellmath__203_0_I10872 (.Y(N12045), .AN(N8271), .B(N8535), .C(N7998));
NAND3XL hyperpropagate_4_1_A_I11464 (.Y(N23383), .A(N9126), .B(N7910), .C(N8779));
NOR2X1 hyperpropagate_4_1_A_I11465 (.Y(N12405), .A(N23383), .B(N8244));
NAND3XL hyperpropagate_4_1_A_I11466 (.Y(N23391), .A(N8675), .B(N8627), .C(N8319));
NOR2X1 hyperpropagate_4_1_A_I11467 (.Y(N12755), .A(N8479), .B(N23391));
NOR4X1 inst_cellmath__203_0_I11221 (.Y(N13112), .A(N8346), .B(N8895), .C(N8455), .D(N7923));
NOR4X1 inst_cellmath__203_0_I11001 (.Y(N11819), .A(N8864), .B(N8655), .C(N8647), .D(N8174));
NOR3BX1 inst_cellmath__203_0_I10878 (.Y(N12192), .AN(N9085), .B(N8887), .C(N8352));
NAND3XL hyperpropagate_4_1_A_I11468 (.Y(N23399), .A(N8815), .B(N8986), .C(N7950));
NOR2X1 hyperpropagate_4_1_A_I11469 (.Y(N12559), .A(N8124), .B(N23399));
INVX1 inst_cellmath__203_0_I3245 (.Y(N12893), .A(inst_cellmath__197[16]));
NAND3XL hyperpropagate_4_1_A_I11470 (.Y(N23407), .A(N8371), .B(N8808), .C(N8596));
NOR2X1 hyperpropagate_4_1_A_I11471 (.Y(N13273), .A(N8485), .B(N23407));
NOR4BX4 inst_cellmath__203_0_I11222 (.Y(N11979), .AN(N8034), .B(N8835), .C(N8720), .D(N7926));
NAND3XL hyperpropagate_4_1_A_I11472 (.Y(N23415), .A(N9042), .B(N8052), .C(N8695));
NOR2X1 hyperpropagate_4_1_A_I11473 (.Y(N12342), .A(N23415), .B(N8589));
MX2X1 inst_cellmath__203_0_I10745 (.Y(N11910), .A(N10755), .B(N10897), .S0(N10460));
INVX2 inst_cellmath__203_0_I10580 (.Y(N23285), .A(N11910));
INVXL inst_cellmath__203_0_I10585 (.Y(N23290), .A(N23285));
INVXL inst_cellmath__203_0_I10583 (.Y(N23288), .A(N23285));
INVX2 inst_cellmath__203_0_I10581 (.Y(N23286), .A(N23285));
NOR2XL inst_cellmath__203_0_I3251 (.Y(N13299), .A(N23290), .B(N12468));
NOR2XL inst_cellmath__203_0_I3252 (.Y(N12367), .A(N23290), .B(N12807));
NOR2XL inst_cellmath__203_0_I3253 (.Y(N13069), .A(N23290), .B(N13175));
NOR2XL inst_cellmath__203_0_I3254 (.Y(N12154), .A(N23290), .B(N11881));
NOR2XL inst_cellmath__203_0_I3255 (.Y(N12856), .A(N23290), .B(N12253));
NOR2XL inst_cellmath__203_0_I3256 (.Y(N11939), .A(N23288), .B(N12618));
NOR2XL inst_cellmath__203_0_I3257 (.Y(N12665), .A(N23288), .B(N12956));
NOR2XL inst_cellmath__203_0_I3258 (.Y(N11719), .A(N23288), .B(N13340));
NOR2XL inst_cellmath__203_0_I3259 (.Y(N12454), .A(N23288), .B(N12045));
NOR2XL inst_cellmath__203_0_I3260 (.Y(N13161), .A(N23288), .B(N12405));
NOR2XL inst_cellmath__203_0_I3261 (.Y(N12241), .A(N23288), .B(N12755));
NOR2XL inst_cellmath__203_0_I3262 (.Y(N12943), .A(N23288), .B(N13112));
NOR2XL inst_cellmath__203_0_I3263 (.Y(N12032), .A(N23288), .B(N11819));
NOR2XL inst_cellmath__203_0_I3264 (.Y(N12746), .A(N23286), .B(N12192));
NOR2XL inst_cellmath__203_0_I3265 (.Y(N11808), .A(N23286), .B(N12559));
NOR2XL inst_cellmath__203_0_I3266 (.Y(N12545), .A(N11910), .B(N12893));
NOR2XL inst_cellmath__203_0_I3267 (.Y(N13263), .A(N11910), .B(N13273));
NOR2X1 inst_cellmath__203_0_I3268 (.Y(N12332), .A(N11979), .B(N23286));
NOR2XL inst_cellmath__203_0_I3269 (.Y(N13033), .A(N11910), .B(N12342));
INVX1 inst_cellmath__203_0_I3271 (.Y(N13137), .A(inst_cellmath__198[18]));
BUFX2 inst_cellmath__203_0_I10746 (.Y(N23296), .A(N13137));
NAND2BX2 inst_cellmath__203_0_I10747 (.Y(N12725), .AN(inst_cellmath__198[19]), .B(inst_cellmath__198[18]));
INVXL inst_cellmath__203_0_I3273 (.Y(N13073), .A(inst_cellmath__198[19]));
NOR2XL inst_cellmath__203_0_I3274 (.Y(N12077), .A(N12104), .B(N23296));
MXI2XL inst_cellmath__203_0_I3275 (.Y(inst_cellmath__203__W1[1]), .A(N13073), .B(N12725), .S0(N12077));
MXI2XL inst_cellmath__203_0_I3276 (.Y(N12013), .A(N12468), .B(N12104), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3277 (.Y(inst_cellmath__203__W0[2]), .A(N13073), .B(N12725), .S0(N12013));
MXI2XL inst_cellmath__203_0_I3278 (.Y(N11950), .A(N12807), .B(N12468), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3279 (.Y(N12766), .A(N13073), .B(N12725), .S0(N11950));
MXI2XL inst_cellmath__203_0_I3280 (.Y(N11879), .A(N13175), .B(N12807), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3281 (.Y(N13128), .A(N13073), .B(N12725), .S0(N11879));
MXI2XL inst_cellmath__203_0_I3282 (.Y(N11817), .A(N11881), .B(N13175), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3283 (.Y(N11835), .A(N13073), .B(N12725), .S0(N11817));
MXI2XL inst_cellmath__203_0_I3284 (.Y(N11755), .A(N12253), .B(N11881), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3285 (.Y(N12208), .A(N13073), .B(N12725), .S0(N11755));
MXI2XL inst_cellmath__203_0_I3286 (.Y(N11690), .A(N12618), .B(N12253), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3287 (.Y(N12574), .A(N13073), .B(N12725), .S0(N11690));
MXI2XL inst_cellmath__203_0_I3288 (.Y(N13301), .A(N12956), .B(N12618), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3289 (.Y(N12908), .A(N13073), .B(N12725), .S0(N13301));
MXI2XL inst_cellmath__203_0_I3290 (.Y(N13232), .A(N13340), .B(N12956), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3291 (.Y(N13291), .A(N13073), .B(N12725), .S0(N13232));
MXI2XL inst_cellmath__203_0_I3292 (.Y(N13164), .A(N12045), .B(N13340), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3293 (.Y(N11997), .A(N13073), .B(N12725), .S0(N13164));
MXI2XL inst_cellmath__203_0_I3294 (.Y(N13101), .A(N12405), .B(N12045), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3295 (.Y(N12356), .A(N13073), .B(N12725), .S0(N13101));
MXI2XL inst_cellmath__203_0_I3296 (.Y(N13035), .A(N12755), .B(N12405), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3297 (.Y(N12712), .A(N13073), .B(N12725), .S0(N13035));
MXI2XL inst_cellmath__203_0_I3298 (.Y(N12972), .A(N13112), .B(N12755), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3299 (.Y(N13063), .A(N13073), .B(N12725), .S0(N12972));
MXI2XL inst_cellmath__203_0_I3300 (.Y(N12912), .A(N11819), .B(N13112), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3301 (.Y(N11773), .A(N13073), .B(N12725), .S0(N12912));
MXI2XL inst_cellmath__203_0_I3302 (.Y(N12852), .A(N12192), .B(N11819), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3303 (.Y(N12146), .A(N13073), .B(N12725), .S0(N12852));
MXI2XL inst_cellmath__203_0_I3304 (.Y(N12792), .A(N12559), .B(N12192), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3305 (.Y(N12511), .A(N13073), .B(N12725), .S0(N12792));
MXI2XL inst_cellmath__203_0_I3306 (.Y(N12739), .A(N12893), .B(N12559), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3307 (.Y(N12848), .A(N13073), .B(N12725), .S0(N12739));
MXI2XL inst_cellmath__203_0_I3308 (.Y(N12686), .A(N13273), .B(N12893), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3309 (.Y(N13223), .A(N13073), .B(N12725), .S0(N12686));
MXI2XL inst_cellmath__203_0_I3310 (.Y(N12627), .A(N11979), .B(N13273), .S0(N23296));
MXI2XL inst_cellmath__203_0_I3311 (.Y(N11932), .A(N13073), .B(N12725), .S0(N12627));
MXI2XL inst_cellmath__203_0_I3312 (.Y(N12569), .A(N12342), .B(N11979), .S0(N13137));
MXI2XL inst_cellmath__203_0_I3313 (.Y(N12296), .A(N13073), .B(N12725), .S0(N12569));
NAND2XL inst_cellmath__203_0_I3314 (.Y(N12506), .A(N12342), .B(N13137));
MXI2XL inst_cellmath__203_0_I3315 (.Y(N12659), .A(N13073), .B(N12725), .S0(N12506));
OR2XL inst_cellmath__203_0_I3317 (.Y(N13149), .A(inst_cellmath__198[19]), .B(inst_cellmath__198[20]));
AOI21XL inst_cellmath__203_0_I10636 (.Y(N13156), .A0(inst_cellmath__198[20]), .A1(inst_cellmath__198[19]), .B0(inst_cellmath__198[21]));
CLKXOR2X1 inst_cellmath__203_0_I3319 (.Y(N12521), .A(inst_cellmath__198[20]), .B(inst_cellmath__198[19]));
INVX3 inst_cellmath__203_0_I3320 (.Y(N12309), .A(N12521));
NAND2X1 inst_cellmath__203_0_I3321 (.Y(N12244), .A(inst_cellmath__198[21]), .B(N13149));
INVXL inst_cellmath__203_0_I3322 (.Y(N12609), .A(N13156));
NOR2XL inst_cellmath__203_0_I3323 (.Y(N12166), .A(N12104), .B(N12309));
MXI2XL inst_cellmath__203_0_I3324 (.Y(inst_cellmath__203__W0[3]), .A(N12609), .B(N12244), .S0(N12166));
MXI2XL inst_cellmath__203_0_I3325 (.Y(N12108), .A(N12104), .B(N12468), .S0(N12521));
MXI2XL inst_cellmath__203_0_I3326 (.Y(N13322), .A(N12609), .B(N12244), .S0(N12108));
MXI2XL inst_cellmath__203_0_I3327 (.Y(N12048), .A(N12807), .B(N12468), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3328 (.Y(N12024), .A(N12609), .B(N12244), .S0(N12048));
MXI2XL inst_cellmath__203_0_I3329 (.Y(N11981), .A(N13175), .B(N12807), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3330 (.Y(N12385), .A(N12609), .B(N12244), .S0(N11981));
MXI2XL inst_cellmath__203_0_I3331 (.Y(N11914), .A(N11881), .B(N13175), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3332 (.Y(N12736), .A(N12609), .B(N12244), .S0(N11914));
MXI2XL inst_cellmath__203_0_I3333 (.Y(N11847), .A(N12253), .B(N11881), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3334 (.Y(N13094), .A(N12609), .B(N12244), .S0(N11847));
MXI2XL inst_cellmath__203_0_I3335 (.Y(N11788), .A(N12618), .B(N12253), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3336 (.Y(N11801), .A(N12609), .B(N12244), .S0(N11788));
MXI2XL inst_cellmath__203_0_I3337 (.Y(N11724), .A(N12956), .B(N12618), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3338 (.Y(N12172), .A(N12609), .B(N12244), .S0(N11724));
MXI2XL inst_cellmath__203_0_I3339 (.Y(N13336), .A(N13340), .B(N12956), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3340 (.Y(N12538), .A(N12609), .B(N12244), .S0(N13336));
MXI2XL inst_cellmath__203_0_I3341 (.Y(N13269), .A(N12045), .B(N13340), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3342 (.Y(N12875), .A(N12609), .B(N12244), .S0(N13269));
MXI2XL inst_cellmath__203_0_I3343 (.Y(N13201), .A(N12405), .B(N12045), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3344 (.Y(N13255), .A(N12609), .B(N12244), .S0(N13201));
MXI2XL inst_cellmath__203_0_I3345 (.Y(N13134), .A(N12755), .B(N12405), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3346 (.Y(N11961), .A(N12609), .B(N12244), .S0(N13134));
MXI2XL inst_cellmath__203_0_I3347 (.Y(N13070), .A(N13112), .B(N12755), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3348 (.Y(N12325), .A(N12609), .B(N12244), .S0(N13070));
MXI2XL inst_cellmath__203_0_I3349 (.Y(N13005), .A(N11819), .B(N13112), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3350 (.Y(N12685), .A(N12609), .B(N12244), .S0(N13005));
MXI2XL inst_cellmath__203_0_I3351 (.Y(N12944), .A(N12192), .B(N11819), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3352 (.Y(N13026), .A(N12609), .B(N12244), .S0(N12944));
MXI2XL inst_cellmath__203_0_I3353 (.Y(N12881), .A(N12559), .B(N12192), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3354 (.Y(N11739), .A(N12609), .B(N12244), .S0(N12881));
MXI2XL inst_cellmath__203_0_I3355 (.Y(N12822), .A(N12893), .B(N12559), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3356 (.Y(N12116), .A(N12609), .B(N12244), .S0(N12822));
MXI2XL inst_cellmath__203_0_I3357 (.Y(N12767), .A(N13273), .B(N12893), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3358 (.Y(N12475), .A(N12609), .B(N12244), .S0(N12767));
MXI2XL inst_cellmath__203_0_I3359 (.Y(N12713), .A(N11979), .B(N13273), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3360 (.Y(N12817), .A(N12609), .B(N12244), .S0(N12713));
MXI2XL inst_cellmath__203_0_I3361 (.Y(N12660), .A(N12342), .B(N11979), .S0(N12309));
MXI2XL inst_cellmath__203_0_I3362 (.Y(N13187), .A(N12609), .B(N12244), .S0(N12660));
NAND2XL inst_cellmath__203_0_I3363 (.Y(N12600), .A(N12342), .B(N12309));
MXI2XL inst_cellmath__203_0_I3364 (.Y(N11892), .A(N12609), .B(N12244), .S0(N12600));
NAND2XL inst_cellmath__203_0_I3366 (.Y(N13252), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
NOR2XL andori2bb1_A_I11474 (.Y(N23421), .A(inst_cellmath__198[22]), .B(inst_cellmath__198[21]));
NOR2XL andori2bb1_A_I11475 (.Y(N12410), .A(N23421), .B(N23282));
CLKXOR2X1 inst_cellmath__203_0_I3368 (.Y(N12036), .A(inst_cellmath__198[21]), .B(inst_cellmath__198[22]));
INVX3 inst_cellmath__203_0_I3369 (.Y(N12184), .A(N12036));
NAND2X2 inst_cellmath__203_0_I3370 (.Y(N12125), .A(N13252), .B(N23282));
INVX1 inst_cellmath__203_0_I3371 (.Y(N12486), .A(N12410));
NOR2XL inst_cellmath__203_0_I3372 (.Y(N12262), .A(N12104), .B(N12184));
MXI2XL inst_cellmath__203_0_I3373 (.Y(N12198), .A(N12486), .B(N12125), .S0(N12262));
MXI2XL inst_cellmath__203_0_I3374 (.Y(N12199), .A(N12104), .B(N12468), .S0(N12036));
MXI2XL inst_cellmath__203_0_I3375 (.Y(N12568), .A(N12486), .B(N12125), .S0(N12199));
MXI2XL inst_cellmath__203_0_I3376 (.Y(N12138), .A(N12807), .B(N12468), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3377 (.Y(N12901), .A(N12486), .B(N12125), .S0(N12138));
MXI2XL inst_cellmath__203_0_I3378 (.Y(N12080), .A(N13175), .B(N12807), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3379 (.Y(N13282), .A(N12486), .B(N12125), .S0(N12080));
MXI2XL inst_cellmath__203_0_I3380 (.Y(N12014), .A(N11881), .B(N13175), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3381 (.Y(N11988), .A(N12486), .B(N12125), .S0(N12014));
MXI2XL inst_cellmath__203_0_I3382 (.Y(N11952), .A(N12253), .B(N11881), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3383 (.Y(N12348), .A(N12486), .B(N12125), .S0(N11952));
MXI2XL inst_cellmath__203_0_I3384 (.Y(N11884), .A(N12618), .B(N12253), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3385 (.Y(N12705), .A(N12486), .B(N12125), .S0(N11884));
MXI2XL inst_cellmath__203_0_I3386 (.Y(N11820), .A(N12956), .B(N12618), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3387 (.Y(N13056), .A(N12486), .B(N12125), .S0(N11820));
MXI2XL inst_cellmath__203_0_I3388 (.Y(N11758), .A(N13340), .B(N12956), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3389 (.Y(N11764), .A(N12486), .B(N12125), .S0(N11758));
MXI2XL inst_cellmath__203_0_I3390 (.Y(N11693), .A(N12045), .B(N13340), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3391 (.Y(N12137), .A(N12486), .B(N12125), .S0(N11693));
MXI2XL inst_cellmath__203_0_I3392 (.Y(N13303), .A(N12405), .B(N12045), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3393 (.Y(N12504), .A(N12486), .B(N12125), .S0(N13303));
MXI2XL inst_cellmath__203_0_I3394 (.Y(N13234), .A(N12755), .B(N12405), .S0(N12184));
MXI2X1 inst_cellmath__203_0_I3395 (.Y(N12841), .A(N12486), .B(N12125), .S0(N13234));
MXI2XL inst_cellmath__203_0_I3396 (.Y(N13167), .A(N13112), .B(N12755), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3397 (.Y(N13214), .A(N12486), .B(N12125), .S0(N13167));
MXI2XL inst_cellmath__203_0_I3398 (.Y(N13104), .A(N11819), .B(N13112), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3399 (.Y(N11922), .A(N12486), .B(N12125), .S0(N13104));
MXI2XL inst_cellmath__203_0_I3400 (.Y(N13037), .A(N12192), .B(N11819), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3401 (.Y(N12288), .A(N12486), .B(N12125), .S0(N13037));
MXI2XL inst_cellmath__203_0_I3402 (.Y(N12976), .A(N12559), .B(N12192), .S0(N12184));
MXI2X1 inst_cellmath__203_0_I3403 (.Y(N12652), .A(N12486), .B(N12125), .S0(N12976));
MXI2XL inst_cellmath__203_0_I3404 (.Y(N12915), .A(N12893), .B(N12559), .S0(N12184));
MXI2X1 inst_cellmath__203_0_I3405 (.Y(N12993), .A(N12486), .B(N12125), .S0(N12915));
MXI2XL inst_cellmath__203_0_I3406 (.Y(N12855), .A(N13273), .B(N12893), .S0(N12184));
MXI2X1 inst_cellmath__203_0_I3407 (.Y(N11701), .A(N12486), .B(N12125), .S0(N12855));
MXI2XL inst_cellmath__203_0_I3408 (.Y(N12795), .A(N11979), .B(N13273), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3409 (.Y(N12079), .A(N12486), .B(N12125), .S0(N12795));
MXI2XL inst_cellmath__203_0_I3410 (.Y(N12743), .A(N12342), .B(N11979), .S0(N12184));
MXI2XL inst_cellmath__203_0_I3411 (.Y(N12440), .A(N12486), .B(N12125), .S0(N12743));
NAND2XL inst_cellmath__203_0_I3412 (.Y(N12690), .A(N12342), .B(N12184));
MXI2XL inst_cellmath__203_0_I3413 (.Y(N12784), .A(N12486), .B(N12125), .S0(N12690));
NAND2XL inst_cellmath__203_0_I3415 (.Y(N11683), .A(inst_cellmath__198[24]), .B(N23282));
NAND2BXL inst_cellmath__203_0_I29536 (.Y(N45195), .AN(N10552), .B(N10682));
XNOR2X1 inst_cellmath__203_0_I29663 (.Y(N45518), .A(N45195), .B(N10899));
XNOR2X1 inst_cellmath__203_0_I29664 (.Y(N45533), .A(N45195), .B(N10400));
MX2X1 inst_cellmath__203_0_I29666 (.Y(inst_cellmath__198[25]), .A(N45518), .B(N45533), .S0(N10407));
NOR2XL andori2bb1_A_I30587 (.Y(N45799), .A(N23282), .B(inst_cellmath__198[24]));
NOR2XL andori2bb1_A_I30588 (.Y(N13312), .A(N45799), .B(inst_cellmath__198[25]));
CLKXOR2X1 inst_cellmath__203_0_I3417 (.Y(N12826), .A(inst_cellmath__198[23]), .B(inst_cellmath__198[24]));
CLKINVX4 inst_cellmath__203_0_I3418 (.Y(N12974), .A(N12826));
AND2XL inst_cellmath__203_0_I10406 (.Y(N23226), .A(N11683), .B(inst_cellmath__198[25]));
INVX2 inst_cellmath__203_0_I10407 (.Y(N12577), .A(N23226));
INVX2 inst_cellmath__203_0_I3421 (.Y(N12914), .A(N13312));
NOR2XL inst_cellmath__203_0_I3422 (.Y(N12354), .A(N12104), .B(N12974));
MXI2XL inst_cellmath__203_0_I3423 (.Y(N13083), .A(N12914), .B(N12577), .S0(N12354));
MXI2XL inst_cellmath__203_0_I3424 (.Y(N12294), .A(N12468), .B(N12104), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3425 (.Y(N11792), .A(N12914), .B(N12577), .S0(N12294));
MXI2XL inst_cellmath__203_0_I3426 (.Y(N12231), .A(N12807), .B(N12468), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3427 (.Y(N12164), .A(N12914), .B(N12577), .S0(N12231));
MXI2XL inst_cellmath__203_0_I3428 (.Y(N12170), .A(N13175), .B(N12807), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3429 (.Y(N12531), .A(N12914), .B(N12577), .S0(N12170));
MXI2XL inst_cellmath__203_0_I3430 (.Y(N12113), .A(N11881), .B(N13175), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3431 (.Y(N12868), .A(N12914), .B(N12577), .S0(N12113));
MXI2XL inst_cellmath__203_0_I3432 (.Y(N12052), .A(N12253), .B(N11881), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3433 (.Y(N13243), .A(N12914), .B(N12577), .S0(N12052));
MXI2XL inst_cellmath__203_0_I3434 (.Y(N11985), .A(N12618), .B(N12253), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3435 (.Y(N11951), .A(N12914), .B(N12577), .S0(N11985));
MXI2XL inst_cellmath__203_0_I3436 (.Y(N11919), .A(N12956), .B(N12618), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3437 (.Y(N12317), .A(N12914), .B(N12577), .S0(N11919));
MXI2XL inst_cellmath__203_0_I3438 (.Y(N11852), .A(N13340), .B(N12956), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3439 (.Y(N12676), .A(N12914), .B(N12577), .S0(N11852));
MXI2XL inst_cellmath__203_0_I3440 (.Y(N11790), .A(N12045), .B(N13340), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3441 (.Y(N13017), .A(N12914), .B(N12577), .S0(N11790));
MXI2XL inst_cellmath__203_0_I3442 (.Y(N11727), .A(N12405), .B(N12045), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3443 (.Y(N11729), .A(N12914), .B(N12577), .S0(N11727));
MXI2XL inst_cellmath__203_0_I3444 (.Y(N13339), .A(N12755), .B(N12405), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3445 (.Y(N12105), .A(N12914), .B(N12577), .S0(N13339));
MXI2X1 inst_cellmath__203_0_I3446 (.Y(N13272), .A(N13112), .B(N12755), .S0(N12974));
MXI2X1 inst_cellmath__203_0_I3447 (.Y(N12469), .A(N12914), .B(N12577), .S0(N13272));
MXI2XL inst_cellmath__203_0_I3448 (.Y(N13203), .A(N11819), .B(N13112), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3449 (.Y(N12809), .A(N12914), .B(N12577), .S0(N13203));
MXI2XL inst_cellmath__203_0_I3450 (.Y(N13136), .A(N12192), .B(N11819), .S0(N12974));
MXI2X1 inst_cellmath__203_0_I3451 (.Y(N13176), .A(N12914), .B(N12577), .S0(N13136));
MXI2XL inst_cellmath__203_0_I3452 (.Y(N13072), .A(N12559), .B(N12192), .S0(N12974));
MXI2X1 inst_cellmath__203_0_I3453 (.Y(N11883), .A(N12914), .B(N12577), .S0(N13072));
MXI2XL inst_cellmath__203_0_I3454 (.Y(N13007), .A(N12893), .B(N12559), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3455 (.Y(N12255), .A(N12914), .B(N12577), .S0(N13007));
MXI2XL inst_cellmath__203_0_I3456 (.Y(N12947), .A(N13273), .B(N12893), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3457 (.Y(N12619), .A(N12914), .B(N12577), .S0(N12947));
MXI2XL inst_cellmath__203_0_I3458 (.Y(N12885), .A(N11979), .B(N13273), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3459 (.Y(N12958), .A(N12914), .B(N12577), .S0(N12885));
MXI2XL inst_cellmath__203_0_I3460 (.Y(N12824), .A(N12342), .B(N11979), .S0(N12974));
MXI2XL inst_cellmath__203_0_I3461 (.Y(N11668), .A(N12914), .B(N12577), .S0(N12824));
NAND2XL inst_cellmath__203_0_I3462 (.Y(N12769), .A(N12342), .B(N12974));
MXI2XL inst_cellmath__203_0_I3463 (.Y(N12046), .A(N12914), .B(N12577), .S0(N12769));
NAND2BXL inst_cellmath__203_0_I29537 (.Y(N45203), .AN(N10818), .B(N10957));
INVXL inst_cellmath__203_0_I29535 (.Y(N45190), .A(N10652));
NOR2BX1 inst_cellmath__203_0_I29542 (.Y(N45206), .AN(N10777), .B(N45190));
XNOR2X1 inst_cellmath__203_0_I29667 (.Y(N45526), .A(N45203), .B(N45190));
XOR2XL inst_cellmath__203_0_I29668 (.Y(N45530), .A(N45203), .B(N45206));
MX2X1 inst_cellmath__203_0_I29669 (.Y(inst_cellmath__198[26]), .A(N45526), .B(N45530), .S0(N10407));
NOR2XL inst_cellmath__203_0_I3464 (.Y(N12716), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NAND2XL inst_cellmath__203_0_I3465 (.Y(N11779), .A(inst_cellmath__198[26]), .B(inst_cellmath__198[25]));
NOR2X1 inst_cellmath__203_0_I3466 (.Y(N12562), .A(N12716), .B(inst_cellmath__198[27]));
CLKXOR2X1 inst_cellmath__203_0_I29670 (.Y(N23303), .A(inst_cellmath__198[25]), .B(inst_cellmath__198[26]));
MXI2XL inst_cellmath__203_0_I29671 (.Y(N45525), .A(N45518), .B(N45533), .S0(N10407));
MXI2X1 inst_cellmath__203_0_I29672 (.Y(N12152), .A(inst_cellmath__198[25]), .B(N45525), .S0(inst_cellmath__198[26]));
BUFX3 inst_cellmath__203_0_I11488 (.Y(N23302), .A(N12152));
INVX2 inst_cellmath__203_0_I10599 (.Y(N23304), .A(N23303));
NAND2X2 inst_cellmath__203_0_I3470 (.Y(N11715), .A(N11779), .B(inst_cellmath__198[27]));
INVX2 inst_cellmath__203_0_I3471 (.Y(N12092), .A(N12562));
NOR2XL inst_cellmath__203_0_I3472 (.Y(N12449), .A(N12104), .B(N23304));
MXI2XL inst_cellmath__203_0_I3473 (.Y(N12343), .A(N12092), .B(N11715), .S0(N12449));
MXI2XL inst_cellmath__203_0_I3474 (.Y(N12388), .A(N12468), .B(N12104), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3475 (.Y(N12700), .A(N12092), .B(N11715), .S0(N12388));
MXI2XL inst_cellmath__203_0_I3476 (.Y(N12327), .A(N12807), .B(N12468), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3477 (.Y(N13047), .A(N12092), .B(N11715), .S0(N12327));
MXI2XL inst_cellmath__203_0_I3478 (.Y(N12266), .A(N13175), .B(N12807), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3479 (.Y(N11757), .A(N12092), .B(N11715), .S0(N12266));
MXI2XL inst_cellmath__203_0_I3480 (.Y(N12201), .A(N11881), .B(N13175), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3481 (.Y(N12133), .A(N12092), .B(N11715), .S0(N12201));
MXI2XL inst_cellmath__203_0_I3482 (.Y(N12140), .A(N12253), .B(N11881), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3483 (.Y(N12496), .A(N12092), .B(N11715), .S0(N12140));
MXI2XL inst_cellmath__203_0_I3484 (.Y(N12082), .A(N12618), .B(N12253), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3485 (.Y(N12833), .A(N12092), .B(N11715), .S0(N12082));
MXI2XL inst_cellmath__203_0_I3486 (.Y(N12017), .A(N12956), .B(N12618), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3487 (.Y(N13205), .A(N12092), .B(N11715), .S0(N12017));
MXI2XL inst_cellmath__203_0_I3488 (.Y(N11956), .A(N13340), .B(N12956), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3489 (.Y(N11912), .A(N12092), .B(N11715), .S0(N11956));
MXI2X1 inst_cellmath__203_0_I3490 (.Y(N11887), .A(N12045), .B(N13340), .S0(N23302));
MXI2X1 inst_cellmath__203_0_I3491 (.Y(N12282), .A(N12092), .B(N11715), .S0(N11887));
MXI2X1 inst_cellmath__203_0_I3492 (.Y(N11823), .A(N12405), .B(N12045), .S0(N23304));
MXI2X1 inst_cellmath__203_0_I3493 (.Y(N12644), .A(N12092), .B(N11715), .S0(N11823));
MXI2X1 inst_cellmath__203_0_I3494 (.Y(N11761), .A(N12755), .B(N12405), .S0(N23302));
MXI2X1 inst_cellmath__203_0_I3495 (.Y(N12983), .A(N12092), .B(N11715), .S0(N11761));
MXI2X1 inst_cellmath__203_0_I3496 (.Y(N11695), .A(N13112), .B(N12755), .S0(N23302));
MXI2X1 inst_cellmath__203_0_I3497 (.Y(N11692), .A(N12092), .B(N11715), .S0(N11695));
MXI2X1 inst_cellmath__203_0_I3498 (.Y(N13308), .A(N11819), .B(N13112), .S0(N23302));
MXI2X1 inst_cellmath__203_0_I3499 (.Y(N12071), .A(N12092), .B(N11715), .S0(N13308));
MXI2XL inst_cellmath__203_0_I3500 (.Y(N13239), .A(N12192), .B(N11819), .S0(N23302));
MXI2XL inst_cellmath__203_0_I3501 (.Y(N12432), .A(N12092), .B(N11715), .S0(N13239));
MXI2XL inst_cellmath__203_0_I3502 (.Y(N13171), .A(N12559), .B(N12192), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3503 (.Y(N12777), .A(N12092), .B(N11715), .S0(N13171));
MXI2XL inst_cellmath__203_0_I3504 (.Y(N13108), .A(N12893), .B(N12559), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3505 (.Y(N13138), .A(N12092), .B(N11715), .S0(N13108));
MXI2XL inst_cellmath__203_0_I3506 (.Y(N13041), .A(N13273), .B(N12893), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3507 (.Y(N11846), .A(N12092), .B(N11715), .S0(N13041));
MXI2XL inst_cellmath__203_0_I3508 (.Y(N12979), .A(N11979), .B(N13273), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3509 (.Y(N12220), .A(N12092), .B(N11715), .S0(N12979));
MXI2XL inst_cellmath__203_0_I3510 (.Y(N12921), .A(N12342), .B(N11979), .S0(N23304));
MXI2XL inst_cellmath__203_0_I3511 (.Y(N12588), .A(N12092), .B(N11715), .S0(N12921));
NAND2XL inst_cellmath__203_0_I3512 (.Y(N12858), .A(N12342), .B(N23304));
MXI2XL inst_cellmath__203_0_I3513 (.Y(N12925), .A(N12092), .B(N11715), .S0(N12858));
NOR2XL inst_cellmath__203_0_I3514 (.Y(N12798), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
NOR2XL inst_cellmath__203_0_I3516 (.Y(N11785), .A(N12798), .B(inst_cellmath__198[29]));
XOR2X1 inst_cellmath__203_0_I3517 (.Y(N12450), .A(inst_cellmath__198[28]), .B(inst_cellmath__198[27]));
INVX3 inst_cellmath__203_0_I3518 (.Y(N12235), .A(N12450));
OAI2BB1X1 inst_cellmath__203_0_I11232 (.Y(N12177), .A0N(inst_cellmath__198[28]), .A1N(inst_cellmath__198[27]), .B0(inst_cellmath__198[29]));
INVX1 inst_cellmath__203_0_I3520 (.Y(N12542), .A(N11785));
NOR2XL inst_cellmath__203_0_I3521 (.Y(N12548), .A(N12104), .B(N12235));
MXI2XL inst_cellmath__203_0_I3522 (.Y(N13233), .A(N12542), .B(N12177), .S0(N12548));
MXI2XL inst_cellmath__203_0_I3523 (.Y(N12483), .A(N12104), .B(N12468), .S0(N12450));
MXI2XL inst_cellmath__203_0_I3524 (.Y(N11942), .A(N12542), .B(N12177), .S0(N12483));
MXI2XL inst_cellmath__203_0_I3525 (.Y(N12419), .A(N12807), .B(N12468), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3526 (.Y(N12311), .A(N12542), .B(N12177), .S0(N12419));
MXI2XL inst_cellmath__203_0_I3527 (.Y(N12359), .A(N13175), .B(N12807), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3528 (.Y(N12669), .A(N12542), .B(N12177), .S0(N12359));
MXI2XL inst_cellmath__203_0_I3529 (.Y(N12299), .A(N11881), .B(N13175), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3530 (.Y(N13008), .A(N12542), .B(N12177), .S0(N12299));
MXI2XL inst_cellmath__203_0_I3531 (.Y(N12233), .A(N12253), .B(N11881), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3532 (.Y(N11722), .A(N12542), .B(N12177), .S0(N12233));
MXI2XL inst_cellmath__203_0_I3533 (.Y(N12173), .A(N12618), .B(N12253), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3534 (.Y(N12099), .A(N12542), .B(N12177), .S0(N12173));
MXI2XL inst_cellmath__203_0_I3535 (.Y(N12117), .A(N12956), .B(N12618), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3536 (.Y(N12461), .A(N12542), .B(N12177), .S0(N12117));
MXI2XL inst_cellmath__203_0_I3537 (.Y(N12054), .A(N13340), .B(N12956), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3538 (.Y(N12802), .A(N12542), .B(N12177), .S0(N12054));
MXI2XL inst_cellmath__203_0_I3539 (.Y(N11989), .A(N12045), .B(N13340), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3540 (.Y(N13166), .A(N12542), .B(N12177), .S0(N11989));
MXI2XL inst_cellmath__203_0_I3541 (.Y(N11923), .A(N12405), .B(N12045), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3542 (.Y(N11872), .A(N12542), .B(N12177), .S0(N11923));
MXI2XL inst_cellmath__203_0_I3543 (.Y(N11855), .A(N12755), .B(N12405), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3544 (.Y(N12248), .A(N12542), .B(N12177), .S0(N11855));
MXI2XL inst_cellmath__203_0_I3545 (.Y(N11793), .A(N13112), .B(N12755), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3546 (.Y(N12610), .A(N12542), .B(N12177), .S0(N11793));
MXI2XL inst_cellmath__203_0_I3547 (.Y(N11730), .A(N11819), .B(N13112), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3548 (.Y(N12948), .A(N12542), .B(N12177), .S0(N11730));
MXI2XL inst_cellmath__203_0_I3549 (.Y(N11669), .A(N12192), .B(N11819), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3550 (.Y(N13333), .A(N12542), .B(N12177), .S0(N11669));
MXI2XL inst_cellmath__203_0_I3551 (.Y(N13274), .A(N12559), .B(N12192), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3552 (.Y(N12037), .A(N12542), .B(N12177), .S0(N13274));
MXI2XL inst_cellmath__203_0_I3553 (.Y(N13206), .A(N12893), .B(N12559), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3554 (.Y(N12397), .A(N12542), .B(N12177), .S0(N13206));
MXI2XL inst_cellmath__203_0_I3555 (.Y(N13139), .A(N13273), .B(N12893), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3556 (.Y(N12749), .A(N12542), .B(N12177), .S0(N13139));
MXI2XL inst_cellmath__203_0_I3557 (.Y(N13075), .A(N11979), .B(N13273), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3558 (.Y(N13103), .A(N12542), .B(N12177), .S0(N13075));
MXI2XL inst_cellmath__203_0_I3559 (.Y(N13009), .A(N12342), .B(N11979), .S0(N12235));
MXI2XL inst_cellmath__203_0_I3560 (.Y(N11812), .A(N12542), .B(N12177), .S0(N13009));
NAND2XL inst_cellmath__203_0_I3561 (.Y(N12949), .A(N12342), .B(N12235));
MXI2XL inst_cellmath__203_0_I3562 (.Y(N12188), .A(N12542), .B(N12177), .S0(N12949));
OA21X1 inst_cellmath__203_0_I11233 (.Y(N12695), .A0(inst_cellmath__198[30]), .A1(inst_cellmath__198[29]), .B0(inst_cellmath__198[31]));
XNOR2X1 inst_cellmath__203_0_I11234 (.Y(N11744), .A(inst_cellmath__198[30]), .B(inst_cellmath__198[29]));
INVXL inst_cellmath__203_0_I10602 (.Y(N23307), .A(N11744));
INVX2 inst_cellmath__203_0_I10603 (.Y(N23308), .A(N23307));
INVX1 inst_cellmath__203_0_I10604 (.Y(N23309), .A(N11744));
INVX1 inst_cellmath__203_0_I10608 (.Y(N23313), .A(N23309));
INVX2 inst_cellmath__203_0_I10607 (.Y(N23312), .A(N23309));
AO21XL inst_cellmath__203_0_I11236 (.Y(N12968), .A0(inst_cellmath__198[29]), .A1(inst_cellmath__198[30]), .B0(inst_cellmath__198[31]));
INVX1 inst_cellmath__203_0_I3570 (.Y(N11679), .A(N12695));
NOR2XL inst_cellmath__203_0_I3571 (.Y(N12638), .A(N12104), .B(N23313));
MXI2XL inst_cellmath__203_0_I3572 (.Y(N12487), .A(N11679), .B(N12968), .S0(N12638));
MXI2XL inst_cellmath__203_0_I3573 (.Y(N12580), .A(N12468), .B(N12104), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3574 (.Y(N12828), .A(N11679), .B(N12968), .S0(N12580));
MXI2XL inst_cellmath__203_0_I3575 (.Y(N12515), .A(N12807), .B(N12468), .S0(N23313));
MXI2XL inst_cellmath__203_0_I3576 (.Y(N13198), .A(N11679), .B(N12968), .S0(N12515));
MXI2XL inst_cellmath__203_0_I3577 (.Y(N12452), .A(N13175), .B(N12807), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3578 (.Y(N11904), .A(N11679), .B(N12968), .S0(N12452));
MXI2XL inst_cellmath__203_0_I3579 (.Y(N12390), .A(N11881), .B(N13175), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3580 (.Y(N12274), .A(N11679), .B(N12968), .S0(N12390));
MXI2XL inst_cellmath__203_0_I3581 (.Y(N12330), .A(N12253), .B(N11881), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3582 (.Y(N12637), .A(N11679), .B(N12968), .S0(N12330));
MXI2XL inst_cellmath__203_0_I3583 (.Y(N12267), .A(N12618), .B(N12253), .S0(N23308));
MXI2X1 inst_cellmath__203_0_I3584 (.Y(N12975), .A(N11679), .B(N12968), .S0(N12267));
MXI2XL inst_cellmath__203_0_I3585 (.Y(N12206), .A(N12956), .B(N12618), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3586 (.Y(N11687), .A(N11679), .B(N12968), .S0(N12206));
MXI2XL inst_cellmath__203_0_I3587 (.Y(N12144), .A(N13340), .B(N12956), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3588 (.Y(N12068), .A(N11679), .B(N12968), .S0(N12144));
MXI2XL inst_cellmath__203_0_I3589 (.Y(N12086), .A(N12045), .B(N13340), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3590 (.Y(N12424), .A(N11679), .B(N12968), .S0(N12086));
MXI2XL inst_cellmath__203_0_I3591 (.Y(N12022), .A(N12405), .B(N12045), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3592 (.Y(N12771), .A(N11679), .B(N12968), .S0(N12022));
MXI2XL inst_cellmath__203_0_I3593 (.Y(N11960), .A(N12755), .B(N12405), .S0(N23312));
MXI2XL inst_cellmath__203_0_I3594 (.Y(N13132), .A(N11679), .B(N12968), .S0(N11960));
MXI2XL inst_cellmath__203_0_I3595 (.Y(N11891), .A(N13112), .B(N12755), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3596 (.Y(N11841), .A(N11679), .B(N12968), .S0(N11891));
MXI2XL inst_cellmath__203_0_I3597 (.Y(N11827), .A(N11819), .B(N13112), .S0(N23313));
MXI2XL inst_cellmath__203_0_I3598 (.Y(N12213), .A(N11679), .B(N12968), .S0(N11827));
MXI2XL inst_cellmath__203_0_I3599 (.Y(N11763), .A(N12192), .B(N11819), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3600 (.Y(N12579), .A(N11679), .B(N12968), .S0(N11763));
MXI2XL inst_cellmath__203_0_I3601 (.Y(N11700), .A(N12559), .B(N12192), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3602 (.Y(N12918), .A(N11679), .B(N12968), .S0(N11700));
MXI2XL inst_cellmath__203_0_I3603 (.Y(N13311), .A(N12893), .B(N12559), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3604 (.Y(N13295), .A(N11679), .B(N12968), .S0(N13311));
MXI2XL inst_cellmath__203_0_I3605 (.Y(N13242), .A(N13273), .B(N12893), .S0(N23308));
MXI2XL inst_cellmath__203_0_I3606 (.Y(N12004), .A(N11679), .B(N12968), .S0(N13242));
MXI2XL inst_cellmath__203_0_I3607 (.Y(N13174), .A(N11979), .B(N13273), .S0(N23313));
MXI2XL inst_cellmath__203_0_I3608 (.Y(N12365), .A(N11679), .B(N12968), .S0(N13174));
MXI2XL inst_cellmath__203_0_I3609 (.Y(N13111), .A(N12342), .B(N11979), .S0(N23313));
MXI2XL inst_cellmath__203_0_I3610 (.Y(N12718), .A(N11679), .B(N12968), .S0(N13111));
NAND2XL inst_cellmath__203_0_I3611 (.Y(N13045), .A(N12342), .B(N23313));
MXI2XL inst_cellmath__203_0_I3612 (.Y(N13067), .A(N11679), .B(N12968), .S0(N13045));
ADDHX1 inst_cellmath__203_0_I3613 (.CO(N13228), .S(N12514), .A(inst_cellmath__198[31]), .B(inst_cellmath__198[32]));
INVX2 inst_cellmath__203_0_I3614 (.Y(N12058), .A(N12514));
INVX2 inst_cellmath__203_0_I10609 (.Y(N23314), .A(N12058));
CLKINVX6 inst_cellmath__203_0_I10610 (.Y(N23315), .A(N23314));
INVX2 inst_cellmath__203_0_I3615 (.Y(N12414), .A(N13228));
NOR2XL inst_cellmath__203_0_I3616 (.Y(N13159), .A(N23315), .B(N12104));
OAI22XL inst_cellmath__203_0_I3617 (.Y(N12237), .A0(N12104), .A1(N12414), .B0(N23315), .B1(N12468));
OAI22XL inst_cellmath__203_0_I3618 (.Y(N12941), .A0(N12468), .A1(N12414), .B0(N12807), .B1(N23315));
OAI22X1 inst_cellmath__203_0_I3619 (.Y(N12029), .A0(N12807), .A1(N12414), .B0(N23315), .B1(N13175));
OAI22XL inst_cellmath__203_0_I3620 (.Y(N12742), .A0(N13175), .A1(N12414), .B0(N11881), .B1(N23315));
OAI22X1 inst_cellmath__203_0_I3621 (.Y(N11806), .A0(N11881), .A1(N12414), .B0(N23315), .B1(N12253));
OAI22XL inst_cellmath__203_0_I3622 (.Y(N12543), .A0(N12253), .A1(N12414), .B0(N23315), .B1(N12618));
OAI22X1 inst_cellmath__203_0_I3623 (.Y(N13260), .A0(N12618), .A1(N12414), .B0(N23315), .B1(N12956));
OAI22X1 inst_cellmath__203_0_I3624 (.Y(N12329), .A0(N12956), .A1(N12414), .B0(N23315), .B1(N13340));
OAI22XL inst_cellmath__203_0_I3625 (.Y(N13031), .A0(N12414), .A1(N13340), .B0(N12045), .B1(N12058));
OAI22XL inst_cellmath__203_0_I3626 (.Y(N12121), .A0(N12045), .A1(N12414), .B0(N23315), .B1(N12405));
OAI22XL inst_cellmath__203_0_I3627 (.Y(N12821), .A0(N12405), .A1(N12414), .B0(N23315), .B1(N12755));
OAI22XL inst_cellmath__203_0_I3628 (.Y(N11898), .A0(N12755), .A1(N12414), .B0(N23315), .B1(N13112));
OAI22XL inst_cellmath__203_0_I3629 (.Y(N12630), .A0(N13112), .A1(N12414), .B0(N23315), .B1(N11819));
OAI22XL inst_cellmath__203_0_I3630 (.Y(N11682), .A0(N11819), .A1(N12414), .B0(N23315), .B1(N12192));
OAI22XL inst_cellmath__203_0_I3631 (.Y(N12415), .A0(N12192), .A1(N12414), .B0(N23315), .B1(N12559));
OAI22XL inst_cellmath__203_0_I3632 (.Y(N13125), .A0(N12559), .A1(N12414), .B0(N23315), .B1(N12893));
OAI22XL inst_cellmath__203_0_I3633 (.Y(N12205), .A0(N12893), .A1(N12414), .B0(N23315), .B1(N13273));
OAI22XL inst_cellmath__203_0_I3634 (.Y(N12906), .A0(N13273), .A1(N12414), .B0(N23315), .B1(N11979));
OAI22XL inst_cellmath__203_0_I3635 (.Y(N11994), .A0(N11979), .A1(N12414), .B0(N23315), .B1(N12342));
OAI21XL inst_cellmath__203_0_I3636 (.Y(N12710), .A0(N12414), .A1(N12342), .B0(N23315));
AND2XL inst_cellmath__203_0_I3637 (.Y(N13204), .A(N12414), .B(N23315));
AND2X1 inst_cellmath__203_0_I10764 (.Y(N12763), .A(N8033), .B(N9019));
AND2X1 inst_cellmath__203_0_I10765 (.Y(N13123), .A(N8172), .B(N8429));
AND2XL inst_cellmath__203_0_I10766 (.Y(N11832), .A(N9015), .B(N8560));
AND2XL inst_cellmath__203_0_I10767 (.Y(N12203), .A(N8120), .B(N9106));
AND2XL inst_cellmath__203_0_I10768 (.Y(N12570), .A(N8781), .B(N8512));
AND2XL inst_cellmath__203_0_I10769 (.Y(N12905), .A(N8630), .B(N8368));
AND2XL inst_cellmath__203_0_I10770 (.Y(N13287), .A(N8202), .B(N7924));
AND2X1 inst_cellmath__203_0_I10627 (.Y(N11992), .A(N8694), .B(N8175));
AND2XL inst_cellmath__203_0_I10773 (.Y(N12353), .A(N8963), .B(N8665));
AND2XL inst_cellmath__203_0_I10774 (.Y(N12708), .A(N7951), .B(N8932));
AND2XL inst_cellmath__203_0_I10775 (.Y(N13059), .A(N8208), .B(N7932));
INVX1 inst_cellmath__203_0_I3649 (.Y(N11770), .A(N753));
AND2XL inst_cellmath__203_0_I10777 (.Y(N12142), .A(N8108), .B(N9096));
AND3X1 inst_cellmath__203_0_I10778 (.Y(N12507), .A(N8238), .B(N9061), .C(N8200));
AND2X1 inst_cellmath__203_0_I10779 (.Y(N12846), .A(N8173), .B(N8432));
AND4X1 inst_cellmath__203_0_I11264 (.Y(N13218), .A(N7918), .B(N8026), .C(N8711), .D(N8562));
AND2XL inst_cellmath__203_0_I10781 (.Y(N11926), .A(N8638), .B(N8377));
AND2XL inst_cellmath__203_0_I10782 (.Y(N12292), .A(N8905), .B(N8353));
AND2XL inst_cellmath__203_0_I10783 (.Y(N12655), .A(N8597), .B(N8325));
INVXL inst_cellmath__203_0_I3657 (.Y(N12996), .A(N761));
AND2X1 inst_cellmath__203_0_I10785 (.Y(N11707), .A(N8743), .B(N8624));
CLKAND2X2 inst_cellmath__203_0_I10786 (.Y(N12084), .A(N8605), .B(N8345));
INVXL inst_cellmath__203_0_I3660 (.Y(N12443), .A(inst_cellmath__61[0]));
NOR2XL inst_cellmath__203_0_I3661 (.Y(N12602), .A(N12443), .B(N12763));
NOR2XL inst_cellmath__203_0_I3662 (.Y(N13327), .A(N12443), .B(N13123));
NOR2XL inst_cellmath__203_0_I3663 (.Y(N12387), .A(N12443), .B(N11832));
NOR2XL inst_cellmath__203_0_I3664 (.Y(N13096), .A(N12443), .B(N12203));
NOR2XL inst_cellmath__203_0_I3665 (.Y(N12175), .A(N12443), .B(N12570));
NOR2XL inst_cellmath__203_0_I3666 (.Y(N12877), .A(N12443), .B(N12905));
NOR2XL inst_cellmath__203_0_I3667 (.Y(N11965), .A(N12443), .B(N13287));
NOR2XL inst_cellmath__203_0_I3668 (.Y(N12688), .A(N12443), .B(N11992));
NOR2XL inst_cellmath__203_0_I3669 (.Y(N11743), .A(N12443), .B(N12353));
NOR2XL inst_cellmath__203_0_I3670 (.Y(N12478), .A(N12443), .B(N12708));
NOR2XL inst_cellmath__203_0_I3671 (.Y(N13190), .A(N12443), .B(N13059));
NOR2XL inst_cellmath__203_0_I3672 (.Y(N12265), .A(N12443), .B(N11770));
NOR2XL inst_cellmath__203_0_I3673 (.Y(N12966), .A(N12443), .B(N12142));
NOR2XL inst_cellmath__203_0_I3674 (.Y(N12056), .A(N12443), .B(N12507));
NOR2XL inst_cellmath__203_0_I3675 (.Y(N12762), .A(N12443), .B(N12846));
NOR2XL inst_cellmath__203_0_I3676 (.Y(N11830), .A(N12443), .B(N13218));
NOR2XL inst_cellmath__203_0_I3677 (.Y(N12904), .A(N12443), .B(N11926));
NOR2XL inst_cellmath__203_0_I3678 (.Y(N13285), .A(N12443), .B(N12292));
NOR2XL inst_cellmath__203_0_I3679 (.Y(N12352), .A(N12443), .B(N12655));
NOR2XL inst_cellmath__203_0_I3680 (.Y(N11915), .A(N12443), .B(N12996));
NOR2XL inst_cellmath__203_0_I3681 (.Y(N11876), .A(N12443), .B(N11707));
NOR2XL inst_cellmath__203_0_I3682 (.Y(N12845), .A(N12443), .B(N12084));
INVXL inst_cellmath__203_0_I3683 (.Y(N12787), .A(inst_cellmath__61[1]));
OR2XL inst_cellmath__203_0_I3684 (.Y(N13089), .A(N12787), .B(inst_cellmath__61[2]));
NOR2XL inst_cellmath__203_0_I3686 (.Y(N12724), .A(N12763), .B(N12787));
MXI2XL inst_cellmath__203_0_I3687 (.Y(N13148), .A(N10622), .B(N13089), .S0(N12724));
MXI2XL inst_cellmath__203_0_I3688 (.Y(N12668), .A(N13123), .B(N12763), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3689 (.Y(N11857), .A(N10622), .B(N13089), .S0(N12668));
MXI2XL inst_cellmath__203_0_I3690 (.Y(N12608), .A(N11832), .B(N13123), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3691 (.Y(N12227), .A(N10622), .B(N13089), .S0(N12608));
MXI2XL inst_cellmath__203_0_I3692 (.Y(N12550), .A(N12203), .B(N11832), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3693 (.Y(N12595), .A(N10622), .B(N13089), .S0(N12550));
MXI2XL inst_cellmath__203_0_I3694 (.Y(N12485), .A(N12570), .B(N12203), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3695 (.Y(N12934), .A(N10622), .B(N13089), .S0(N12485));
MXI2XL inst_cellmath__203_0_I3696 (.Y(N12421), .A(N12905), .B(N12570), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3697 (.Y(N13316), .A(N10622), .B(N13089), .S0(N12421));
MXI2XL inst_cellmath__203_0_I3698 (.Y(N12362), .A(N13287), .B(N12905), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3699 (.Y(N12016), .A(N10622), .B(N13089), .S0(N12362));
MXI2XL inst_cellmath__203_0_I3700 (.Y(N12303), .A(N11992), .B(N13287), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3701 (.Y(N12380), .A(N10622), .B(N13089), .S0(N12303));
MXI2XL inst_cellmath__203_0_I3702 (.Y(N12234), .A(N12353), .B(N11992), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3703 (.Y(N12732), .A(N10622), .B(N13089), .S0(N12234));
MXI2XL inst_cellmath__203_0_I3704 (.Y(N12176), .A(N12708), .B(N12353), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3705 (.Y(N13086), .A(N10622), .B(N13089), .S0(N12176));
MXI2XL inst_cellmath__203_0_I3706 (.Y(N12119), .A(N13059), .B(N12708), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3707 (.Y(N11794), .A(N10622), .B(N13089), .S0(N12119));
MXI2XL inst_cellmath__203_0_I3708 (.Y(N12057), .A(N11770), .B(N13059), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3709 (.Y(N12167), .A(N10622), .B(N13089), .S0(N12057));
MXI2XL inst_cellmath__203_0_I3710 (.Y(N11991), .A(N12142), .B(N11770), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3711 (.Y(N12533), .A(N10622), .B(N13089), .S0(N11991));
MXI2XL inst_cellmath__203_0_I3712 (.Y(N11925), .A(N12507), .B(N12142), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3713 (.Y(N12871), .A(N10622), .B(N13089), .S0(N11925));
MXI2XL inst_cellmath__203_0_I3714 (.Y(N11858), .A(N12846), .B(N12507), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3715 (.Y(N13248), .A(N10622), .B(N13089), .S0(N11858));
MXI2XL inst_cellmath__203_0_I3716 (.Y(N11795), .A(N13218), .B(N12846), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3717 (.Y(N11954), .A(N10622), .B(N13089), .S0(N11795));
MXI2XL inst_cellmath__203_0_I3718 (.Y(N11734), .A(N11926), .B(N13218), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3719 (.Y(N12319), .A(N10622), .B(N13089), .S0(N11734));
MXI2XL inst_cellmath__203_0_I3720 (.Y(N11672), .A(N12292), .B(N11926), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3721 (.Y(N12680), .A(N10622), .B(N13089), .S0(N11672));
MXI2XL inst_cellmath__203_0_I3722 (.Y(N13278), .A(N12655), .B(N12292), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3723 (.Y(N13020), .A(N10622), .B(N13089), .S0(N13278));
MXI2XL inst_cellmath__203_0_I3724 (.Y(N13209), .A(N12996), .B(N12655), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3725 (.Y(N11732), .A(N10622), .B(N13089), .S0(N13209));
MXI2XL inst_cellmath__203_0_I3726 (.Y(N13141), .A(N11707), .B(N12996), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3727 (.Y(N12110), .A(N10622), .B(N13089), .S0(N13141));
MXI2X1 inst_cellmath__203_0_I3728 (.Y(N13079), .A(N12084), .B(N11707), .S0(N12787));
MXI2XL inst_cellmath__203_0_I3729 (.Y(N12470), .A(N10622), .B(N13089), .S0(N13079));
NOR2BX1 inst_cellmath__203_0_I3730 (.Y(N13013), .AN(N12787), .B(N12084));
MXI2XL inst_cellmath__203_0_I3731 (.Y(N12812), .A(N10622), .B(N13089), .S0(N13013));
XNOR2X1 inst_cellmath__203_0_I10650 (.Y(N23344), .A(inst_cellmath__61[2]), .B(inst_cellmath__61[3]));
NAND2XL inst_cellmath__203_0_I3733 (.Y(N12953), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
NOR2XL inst_cellmath__203_0_I3734 (.Y(N12042), .A(inst_cellmath__61[3]), .B(inst_cellmath__61[2]));
AND2XL inst_cellmath__203_0_I3735 (.Y(N11671), .A(N12953), .B(inst_cellmath__61[4]));
OR2XL inst_cellmath__203_0_I3736 (.Y(N12499), .A(N12042), .B(inst_cellmath__61[4]));
INVXL inst_cellmath__203_0_I3737 (.Y(N12435), .A(N11671));
NOR2XL inst_cellmath__203_0_I3738 (.Y(N12697), .A(N12763), .B(N23344));
MXI2XL inst_cellmath__203_0_I3739 (.Y(N13116), .A(N12435), .B(N12499), .S0(N12697));
MXI2XL inst_cellmath__203_0_I3740 (.Y(N12641), .A(N13123), .B(N12763), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3741 (.Y(N11822), .A(N12435), .B(N12499), .S0(N12641));
MXI2XL inst_cellmath__203_0_I3742 (.Y(N12584), .A(N11832), .B(N13123), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3743 (.Y(N12195), .A(N12435), .B(N12499), .S0(N12584));
MXI2XL inst_cellmath__203_0_I3744 (.Y(N12518), .A(N12203), .B(N11832), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3745 (.Y(N12564), .A(N12435), .B(N12499), .S0(N12518));
MXI2XL inst_cellmath__203_0_I3746 (.Y(N12455), .A(N12570), .B(N12203), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3747 (.Y(N12896), .A(N12435), .B(N12499), .S0(N12455));
MXI2XL inst_cellmath__203_0_I3748 (.Y(N12393), .A(N12905), .B(N12570), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3749 (.Y(N13277), .A(N12435), .B(N12499), .S0(N12393));
MXI2XL inst_cellmath__203_0_I3750 (.Y(N12334), .A(N13287), .B(N12905), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3751 (.Y(N11983), .A(N12435), .B(N12499), .S0(N12334));
MXI2XL inst_cellmath__203_0_I3752 (.Y(N12270), .A(N11992), .B(N13287), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3753 (.Y(N12344), .A(N12435), .B(N12499), .S0(N12270));
MXI2XL inst_cellmath__203_0_I3754 (.Y(N12209), .A(N12353), .B(N11992), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3755 (.Y(N12702), .A(N12435), .B(N12499), .S0(N12209));
MXI2XL inst_cellmath__203_0_I3756 (.Y(N12148), .A(N12708), .B(N12353), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3757 (.Y(N13050), .A(N12435), .B(N12499), .S0(N12148));
MXI2XL inst_cellmath__203_0_I3758 (.Y(N12089), .A(N13059), .B(N12708), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3759 (.Y(N11760), .A(N12435), .B(N12499), .S0(N12089));
MXI2XL inst_cellmath__203_0_I3760 (.Y(N12025), .A(N11770), .B(N13059), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3761 (.Y(N12134), .A(N12435), .B(N12499), .S0(N12025));
MXI2XL inst_cellmath__203_0_I3762 (.Y(N11964), .A(N12142), .B(N11770), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3763 (.Y(N12498), .A(N12435), .B(N12499), .S0(N11964));
MXI2XL inst_cellmath__203_0_I3764 (.Y(N11895), .A(N12507), .B(N12142), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3765 (.Y(N12836), .A(N12435), .B(N12499), .S0(N11895));
MXI2XL inst_cellmath__203_0_I3766 (.Y(N11828), .A(N12846), .B(N12507), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3767 (.Y(N13208), .A(N12435), .B(N12499), .S0(N11828));
MXI2XL inst_cellmath__203_0_I3768 (.Y(N11767), .A(N13218), .B(N12846), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3769 (.Y(N11916), .A(N12435), .B(N12499), .S0(N11767));
MXI2XL inst_cellmath__203_0_I3770 (.Y(N11704), .A(N11926), .B(N13218), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3771 (.Y(N12284), .A(N12435), .B(N12499), .S0(N11704));
MXI2XL inst_cellmath__203_0_I3772 (.Y(N13314), .A(N12292), .B(N11926), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3773 (.Y(N12648), .A(N12435), .B(N12499), .S0(N13314));
MXI2XL inst_cellmath__203_0_I3774 (.Y(N13245), .A(N12655), .B(N12292), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3775 (.Y(N12986), .A(N12435), .B(N12499), .S0(N13245));
MXI2XL inst_cellmath__203_0_I3776 (.Y(N13178), .A(N12996), .B(N12655), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3777 (.Y(N11697), .A(N12435), .B(N12499), .S0(N13178));
MXI2XL inst_cellmath__203_0_I3778 (.Y(N13114), .A(N11707), .B(N12996), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3779 (.Y(N12074), .A(N12435), .B(N12499), .S0(N13114));
MXI2XL inst_cellmath__203_0_I3780 (.Y(N13048), .A(N12084), .B(N11707), .S0(N23344));
MXI2XL inst_cellmath__203_0_I3781 (.Y(N12434), .A(N12435), .B(N12499), .S0(N13048));
NOR2BX1 inst_cellmath__203_0_I10787 (.Y(N12984), .AN(N23344), .B(N12084));
MXI2XL inst_cellmath__203_0_I3783 (.Y(N12780), .A(N12435), .B(N12499), .S0(N12984));
XNOR2X1 inst_cellmath__203_0_I3784 (.Y(N12591), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
NAND2XL inst_cellmath__203_0_I3785 (.Y(N12926), .A(inst_cellmath__61[5]), .B(inst_cellmath__61[4]));
NOR2XL inst_cellmath__203_0_I3786 (.Y(N12009), .A(inst_cellmath__61[4]), .B(inst_cellmath__61[5]));
AND2XL inst_cellmath__203_0_I3787 (.Y(N13307), .A(N12926), .B(N3808));
OR2XL inst_cellmath__203_0_I3788 (.Y(N11946), .A(N12009), .B(N3808));
INVXL inst_cellmath__203_0_I3789 (.Y(N11877), .A(N13307));
NOR2XL inst_cellmath__203_0_I3790 (.Y(N12671), .A(N12763), .B(N12591));
MXI2XL inst_cellmath__203_0_I3791 (.Y(N13077), .A(N11877), .B(N11946), .S0(N12671));
MXI2XL inst_cellmath__203_0_I3792 (.Y(N12612), .A(N13123), .B(N12763), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3793 (.Y(N11787), .A(N11877), .B(N11946), .S0(N12612));
MXI2XL inst_cellmath__203_0_I3794 (.Y(N12553), .A(N11832), .B(N13123), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3795 (.Y(N12162), .A(N11877), .B(N11946), .S0(N12553));
MXI2XL inst_cellmath__203_0_I3796 (.Y(N12489), .A(N12203), .B(N11832), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3797 (.Y(N12526), .A(N11877), .B(N11946), .S0(N12489));
MXI2XL inst_cellmath__203_0_I3798 (.Y(N12425), .A(N12570), .B(N12203), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3799 (.Y(N12862), .A(N11877), .B(N11946), .S0(N12425));
MXI2XL inst_cellmath__203_0_I3800 (.Y(N12366), .A(N12905), .B(N12570), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3801 (.Y(N13238), .A(N11877), .B(N11946), .S0(N12366));
MXI2XL inst_cellmath__203_0_I3802 (.Y(N12305), .A(N13287), .B(N12905), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3803 (.Y(N11944), .A(N11877), .B(N11946), .S0(N12305));
MXI2XL inst_cellmath__203_0_I3804 (.Y(N12238), .A(N11992), .B(N13287), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3805 (.Y(N12313), .A(N11877), .B(N11946), .S0(N12238));
MXI2XL inst_cellmath__203_0_I3806 (.Y(N12179), .A(N12353), .B(N11992), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3807 (.Y(N12673), .A(N11877), .B(N11946), .S0(N12179));
MXI2XL inst_cellmath__203_0_I3808 (.Y(N12122), .A(N12708), .B(N12353), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3809 (.Y(N13011), .A(N11877), .B(N11946), .S0(N12122));
MXI2XL inst_cellmath__203_0_I3810 (.Y(N12060), .A(N13059), .B(N12708), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3811 (.Y(N11723), .A(N11877), .B(N11946), .S0(N12060));
MXI2XL inst_cellmath__203_0_I3812 (.Y(N11995), .A(N11770), .B(N13059), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3813 (.Y(N12101), .A(N11877), .B(N11946), .S0(N11995));
MXI2XL inst_cellmath__203_0_I3814 (.Y(N11929), .A(N12142), .B(N11770), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3815 (.Y(N12463), .A(N11877), .B(N11946), .S0(N11929));
MXI2XL inst_cellmath__203_0_I3816 (.Y(N11862), .A(N12507), .B(N12142), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3817 (.Y(N12804), .A(N11877), .B(N11946), .S0(N11862));
MXI2XL inst_cellmath__203_0_I3818 (.Y(N11799), .A(N12846), .B(N12507), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3819 (.Y(N13170), .A(N11877), .B(N11946), .S0(N11799));
MXI2XL inst_cellmath__203_0_I3820 (.Y(N11737), .A(N13218), .B(N12846), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3821 (.Y(N11875), .A(N11877), .B(N11946), .S0(N11737));
MXI2XL inst_cellmath__203_0_I3822 (.Y(N11675), .A(N11926), .B(N13218), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3823 (.Y(N12250), .A(N11877), .B(N11946), .S0(N11675));
MXI2XL inst_cellmath__203_0_I3824 (.Y(N13280), .A(N12292), .B(N11926), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3825 (.Y(N12614), .A(N11877), .B(N11946), .S0(N13280));
MXI2XL inst_cellmath__203_0_I3826 (.Y(N13212), .A(N12655), .B(N12292), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3827 (.Y(N12951), .A(N11877), .B(N11946), .S0(N13212));
MXI2XL inst_cellmath__203_0_I3828 (.Y(N13145), .A(N12996), .B(N12655), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3829 (.Y(N13335), .A(N11877), .B(N11946), .S0(N13145));
MXI2XL inst_cellmath__203_0_I3830 (.Y(N13082), .A(N11707), .B(N12996), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3831 (.Y(N12041), .A(N11877), .B(N11946), .S0(N13082));
MXI2XL inst_cellmath__203_0_I3832 (.Y(N13016), .A(N12084), .B(N11707), .S0(N12591));
MXI2XL inst_cellmath__203_0_I3833 (.Y(N12399), .A(N11877), .B(N11946), .S0(N13016));
NOR2BX1 inst_cellmath__203_0_I3834 (.Y(N12957), .AN(N12591), .B(N12084));
MXI2XL inst_cellmath__203_0_I3835 (.Y(N12751), .A(N11877), .B(N11946), .S0(N12957));
XNOR2X1 inst_cellmath__203_0_I3836 (.Y(N12555), .A(inst_cellmath__61[7]), .B(N3808));
NAND2XL inst_cellmath__203_0_I3837 (.Y(N12892), .A(inst_cellmath__61[7]), .B(N3808));
NOR2XL inst_cellmath__203_0_I3838 (.Y(N11978), .A(N3808), .B(inst_cellmath__61[7]));
AND2XL inst_cellmath__203_0_I3839 (.Y(N13268), .A(N12892), .B(inst_cellmath__61[8]));
OR2XL inst_cellmath__203_0_I3840 (.Y(N13042), .A(N11978), .B(inst_cellmath__61[8]));
INVXL inst_cellmath__203_0_I3841 (.Y(N12980), .A(N13268));
NOR2XL inst_cellmath__203_0_I3842 (.Y(N12643), .A(N12763), .B(N12555));
MXI2XL inst_cellmath__203_0_I3843 (.Y(N13040), .A(N12980), .B(N13042), .S0(N12643));
MXI2XL inst_cellmath__203_0_I3844 (.Y(N12586), .A(N13123), .B(N12763), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3845 (.Y(N11752), .A(N12980), .B(N13042), .S0(N12586));
MXI2XL inst_cellmath__203_0_I3846 (.Y(N12522), .A(N11832), .B(N13123), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3847 (.Y(N12130), .A(N12980), .B(N13042), .S0(N12522));
MXI2XL inst_cellmath__203_0_I3848 (.Y(N12459), .A(N12203), .B(N11832), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3849 (.Y(N12491), .A(N12980), .B(N13042), .S0(N12459));
MXI2XL inst_cellmath__203_0_I3850 (.Y(N12395), .A(N12570), .B(N12203), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3851 (.Y(N12829), .A(N12980), .B(N13042), .S0(N12395));
MXI2XL inst_cellmath__203_0_I3852 (.Y(N12336), .A(N12905), .B(N12570), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3853 (.Y(N13200), .A(N12980), .B(N13042), .S0(N12336));
MXI2XL inst_cellmath__203_0_I3854 (.Y(N12272), .A(N13287), .B(N12905), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3855 (.Y(N11908), .A(N12980), .B(N13042), .S0(N12272));
MXI2XL inst_cellmath__203_0_I3856 (.Y(N12212), .A(N11992), .B(N13287), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3857 (.Y(N12277), .A(N12980), .B(N13042), .S0(N12212));
MXI2XL inst_cellmath__203_0_I3858 (.Y(N12151), .A(N12353), .B(N11992), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3859 (.Y(N12640), .A(N12980), .B(N13042), .S0(N12151));
MXI2XL inst_cellmath__203_0_I3860 (.Y(N12091), .A(N12708), .B(N12353), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3861 (.Y(N12978), .A(N12980), .B(N13042), .S0(N12091));
MXI2XL inst_cellmath__203_0_I3862 (.Y(N12028), .A(N13059), .B(N12708), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3863 (.Y(N11689), .A(N12980), .B(N13042), .S0(N12028));
MXI2XL inst_cellmath__203_0_I3864 (.Y(N11967), .A(N11770), .B(N13059), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3865 (.Y(N12069), .A(N12980), .B(N13042), .S0(N11967));
MXI2XL inst_cellmath__203_0_I3866 (.Y(N11897), .A(N12142), .B(N11770), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3867 (.Y(N12427), .A(N12980), .B(N13042), .S0(N11897));
MXI2XL inst_cellmath__203_0_I3868 (.Y(N11831), .A(N12507), .B(N12142), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3869 (.Y(N12774), .A(N12980), .B(N13042), .S0(N11831));
MXI2XL inst_cellmath__203_0_I3870 (.Y(N11769), .A(N12846), .B(N12507), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3871 (.Y(N13133), .A(N12980), .B(N13042), .S0(N11769));
MXI2XL inst_cellmath__203_0_I3872 (.Y(N11706), .A(N13218), .B(N12846), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3873 (.Y(N11842), .A(N12980), .B(N13042), .S0(N11706));
MXI2XL inst_cellmath__203_0_I3874 (.Y(N13317), .A(N11926), .B(N13218), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3875 (.Y(N12216), .A(N12980), .B(N13042), .S0(N13317));
MXI2XL inst_cellmath__203_0_I3876 (.Y(N13249), .A(N12292), .B(N11926), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3877 (.Y(N12583), .A(N12980), .B(N13042), .S0(N13249));
MXI2XL inst_cellmath__203_0_I3878 (.Y(N13181), .A(N12655), .B(N12292), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3879 (.Y(N12920), .A(N12980), .B(N13042), .S0(N13181));
MXI2XL inst_cellmath__203_0_I3880 (.Y(N13117), .A(N12996), .B(N12655), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3881 (.Y(N13298), .A(N12980), .B(N13042), .S0(N13117));
MXI2XL inst_cellmath__203_0_I3882 (.Y(N13051), .A(N11707), .B(N12996), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3883 (.Y(N12006), .A(N12980), .B(N13042), .S0(N13051));
MXI2XL inst_cellmath__203_0_I3884 (.Y(N12987), .A(N12084), .B(N11707), .S0(N12555));
MXI2XL inst_cellmath__203_0_I3885 (.Y(N12369), .A(N12980), .B(N13042), .S0(N12987));
NOR2BX1 inst_cellmath__203_0_I3886 (.Y(N12928), .AN(N12555), .B(N12084));
MXI2XL inst_cellmath__203_0_I3887 (.Y(N12721), .A(N12980), .B(N13042), .S0(N12928));
XNOR2X1 inst_cellmath__203_0_I3888 (.Y(N12517), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
NAND2XL inst_cellmath__203_0_I3889 (.Y(N12863), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
NOR2XL inst_cellmath__203_0_I3890 (.Y(N11947), .A(inst_cellmath__61[9]), .B(inst_cellmath__61[8]));
AND2XL inst_cellmath__203_0_I3891 (.Y(N13230), .A(N12863), .B(N3810));
OR2XL inst_cellmath__203_0_I3892 (.Y(N12519), .A(N11947), .B(N3810));
INVXL inst_cellmath__203_0_I3893 (.Y(N12457), .A(N13230));
NOR2XL inst_cellmath__203_0_I3894 (.Y(N12615), .A(N12763), .B(N12517));
MXI2XL inst_cellmath__203_0_I3895 (.Y(N13004), .A(N12457), .B(N12519), .S0(N12615));
MXI2XL inst_cellmath__203_0_I3896 (.Y(N12556), .A(N13123), .B(N12763), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3897 (.Y(N11718), .A(N12457), .B(N12519), .S0(N12556));
MXI2XL inst_cellmath__203_0_I3898 (.Y(N12492), .A(N11832), .B(N13123), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3899 (.Y(N12096), .A(N12457), .B(N12519), .S0(N12492));
MXI2XL inst_cellmath__203_0_I3900 (.Y(N12428), .A(N12203), .B(N11832), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3901 (.Y(N12453), .A(N12457), .B(N12519), .S0(N12428));
MXI2XL inst_cellmath__203_0_I3902 (.Y(N12370), .A(N12570), .B(N12203), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3903 (.Y(N12797), .A(N12457), .B(N12519), .S0(N12370));
MXI2XL inst_cellmath__203_0_I3904 (.Y(N12307), .A(N12905), .B(N12570), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3905 (.Y(N13163), .A(N12457), .B(N12519), .S0(N12307));
MXI2XL inst_cellmath__203_0_I3906 (.Y(N12242), .A(N13287), .B(N12905), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3907 (.Y(N11867), .A(N12457), .B(N12519), .S0(N12242));
MXI2XL inst_cellmath__203_0_I3908 (.Y(N12182), .A(N11992), .B(N13287), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3909 (.Y(N12240), .A(N12457), .B(N12519), .S0(N12182));
MXI2XL inst_cellmath__203_0_I3910 (.Y(N12124), .A(N12353), .B(N11992), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3911 (.Y(N12606), .A(N12457), .B(N12519), .S0(N12124));
MXI2XL inst_cellmath__203_0_I3912 (.Y(N12063), .A(N12708), .B(N12353), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3913 (.Y(N12942), .A(N12457), .B(N12519), .S0(N12063));
MXI2XL inst_cellmath__203_0_I3914 (.Y(N11999), .A(N13059), .B(N12708), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3915 (.Y(N13328), .A(N12457), .B(N12519), .S0(N11999));
MXI2XL inst_cellmath__203_0_I3916 (.Y(N11933), .A(N11770), .B(N13059), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3917 (.Y(N12033), .A(N12457), .B(N12519), .S0(N11933));
MXI2XL inst_cellmath__203_0_I3918 (.Y(N11864), .A(N12142), .B(N11770), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3919 (.Y(N12391), .A(N12457), .B(N12519), .S0(N11864));
MXI2XL inst_cellmath__203_0_I3920 (.Y(N11802), .A(N12507), .B(N12142), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3921 (.Y(N12745), .A(N12457), .B(N12519), .S0(N11802));
MXI2XL inst_cellmath__203_0_I3922 (.Y(N11741), .A(N12846), .B(N12507), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3923 (.Y(N13100), .A(N12457), .B(N12519), .S0(N11741));
MXI2XL inst_cellmath__203_0_I3924 (.Y(N11677), .A(N13218), .B(N12846), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3925 (.Y(N11807), .A(N12457), .B(N12519), .S0(N11677));
MXI2XL inst_cellmath__203_0_I3926 (.Y(N13284), .A(N11926), .B(N13218), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3927 (.Y(N12181), .A(N12457), .B(N12519), .S0(N13284));
MXI2XL inst_cellmath__203_0_I3928 (.Y(N13216), .A(N12292), .B(N11926), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3929 (.Y(N12547), .A(N12457), .B(N12519), .S0(N13216));
MXI2XL inst_cellmath__203_0_I3930 (.Y(N13147), .A(N12655), .B(N12292), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3931 (.Y(N12880), .A(N12457), .B(N12519), .S0(N13147));
MXI2XL inst_cellmath__203_0_I3932 (.Y(N13085), .A(N12996), .B(N12655), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3933 (.Y(N13262), .A(N12457), .B(N12519), .S0(N13085));
MXI2XL inst_cellmath__203_0_I3934 (.Y(N13019), .A(N11707), .B(N12996), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3935 (.Y(N11971), .A(N12457), .B(N12519), .S0(N13019));
MXI2XL inst_cellmath__203_0_I3936 (.Y(N12960), .A(N12084), .B(N11707), .S0(N12517));
MXI2XL inst_cellmath__203_0_I3937 (.Y(N12331), .A(N12457), .B(N12519), .S0(N12960));
NOR2BX1 inst_cellmath__203_0_I3938 (.Y(N12895), .AN(N12517), .B(N12084));
MXI2XL inst_cellmath__203_0_I3939 (.Y(N12692), .A(N12457), .B(N12519), .S0(N12895));
XNOR2X1 inst_cellmath__203_0_I3940 (.Y(N12482), .A(inst_cellmath__61[11]), .B(N3810));
NAND2XL inst_cellmath__203_0_I3941 (.Y(N12835), .A(inst_cellmath__61[11]), .B(N3810));
NOR2XL inst_cellmath__203_0_I3942 (.Y(N11913), .A(inst_cellmath__61[11]), .B(N3810));
AND2XL inst_cellmath__203_0_I3943 (.Y(N13193), .A(N12835), .B(inst_cellmath__61[12]));
OR2XL inst_cellmath__203_0_I3944 (.Y(N12883), .A(N11913), .B(inst_cellmath__61[12]));
INVXL inst_cellmath__203_0_I3945 (.Y(N12484), .A(N13193));
NOR2XL inst_cellmath__203_0_I3946 (.Y(N12590), .A(N12763), .B(N12482));
MXI2XL inst_cellmath__203_0_I3947 (.Y(N12971), .A(N12484), .B(N12883), .S0(N12590));
MXI2XL inst_cellmath__203_0_I3948 (.Y(N12525), .A(N13123), .B(N12763), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3949 (.Y(N11684), .A(N12484), .B(N12883), .S0(N12525));
MXI2XL inst_cellmath__203_0_I3950 (.Y(N12462), .A(N11832), .B(N13123), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3951 (.Y(N12062), .A(N12484), .B(N12883), .S0(N12462));
MXI2XL inst_cellmath__203_0_I3952 (.Y(N12398), .A(N12203), .B(N11832), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3953 (.Y(N12418), .A(N12484), .B(N12883), .S0(N12398));
MXI2XL inst_cellmath__203_0_I3954 (.Y(N12338), .A(N12570), .B(N12203), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3955 (.Y(N12765), .A(N12484), .B(N12883), .S0(N12338));
MXI2XL inst_cellmath__203_0_I3956 (.Y(N12276), .A(N12905), .B(N12570), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3957 (.Y(N13127), .A(N12484), .B(N12883), .S0(N12276));
MXI2XL inst_cellmath__203_0_I3958 (.Y(N12215), .A(N13287), .B(N12905), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3959 (.Y(N11836), .A(N12484), .B(N12883), .S0(N12215));
MXI2XL inst_cellmath__203_0_I3960 (.Y(N12153), .A(N11992), .B(N13287), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3961 (.Y(N12207), .A(N12484), .B(N12883), .S0(N12153));
MXI2XL inst_cellmath__203_0_I3962 (.Y(N12094), .A(N12353), .B(N11992), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3963 (.Y(N12573), .A(N12484), .B(N12883), .S0(N12094));
MXI2XL inst_cellmath__203_0_I3964 (.Y(N12031), .A(N12708), .B(N12353), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3965 (.Y(N12910), .A(N12484), .B(N12883), .S0(N12031));
MXI2XL inst_cellmath__203_0_I3966 (.Y(N11969), .A(N13059), .B(N12708), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3967 (.Y(N13290), .A(N12484), .B(N12883), .S0(N11969));
MXI2XL inst_cellmath__203_0_I3968 (.Y(N11899), .A(N11770), .B(N13059), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3969 (.Y(N11996), .A(N12484), .B(N12883), .S0(N11899));
MXI2XL inst_cellmath__203_0_I3970 (.Y(N11834), .A(N12142), .B(N11770), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3971 (.Y(N12358), .A(N12484), .B(N12883), .S0(N11834));
MXI2XL inst_cellmath__203_0_I3972 (.Y(N11772), .A(N12507), .B(N12142), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3973 (.Y(N12711), .A(N12484), .B(N12883), .S0(N11772));
MXI2XL inst_cellmath__203_0_I3974 (.Y(N11710), .A(N12846), .B(N12507), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3975 (.Y(N13062), .A(N12484), .B(N12883), .S0(N11710));
MXI2XL inst_cellmath__203_0_I3976 (.Y(N13321), .A(N13218), .B(N12846), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3977 (.Y(N11775), .A(N12484), .B(N12883), .S0(N13321));
MXI2XL inst_cellmath__203_0_I3978 (.Y(N13251), .A(N11926), .B(N13218), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3979 (.Y(N12145), .A(N12484), .B(N12883), .S0(N13251));
MXI2XL inst_cellmath__203_0_I3980 (.Y(N13184), .A(N12292), .B(N11926), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3981 (.Y(N12510), .A(N12484), .B(N12883), .S0(N13184));
MXI2XL inst_cellmath__203_0_I3982 (.Y(N13120), .A(N12655), .B(N12292), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3983 (.Y(N12850), .A(N12484), .B(N12883), .S0(N13120));
MXI2XL inst_cellmath__203_0_I3984 (.Y(N13053), .A(N12996), .B(N12655), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3985 (.Y(N13222), .A(N12484), .B(N12883), .S0(N13053));
MXI2XL inst_cellmath__203_0_I3986 (.Y(N12990), .A(N11707), .B(N12996), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3987 (.Y(N11931), .A(N12484), .B(N12883), .S0(N12990));
MXI2XL inst_cellmath__203_0_I3988 (.Y(N12931), .A(N12084), .B(N11707), .S0(N12482));
MXI2XL inst_cellmath__203_0_I3989 (.Y(N12298), .A(N12484), .B(N12883), .S0(N12931));
NOR2BX1 inst_cellmath__203_0_I3990 (.Y(N12866), .AN(N12482), .B(N12084));
MXI2XL inst_cellmath__203_0_I3991 (.Y(N12658), .A(N12484), .B(N12883), .S0(N12866));
XNOR2X1 inst_cellmath__203_0_I3992 (.Y(N12448), .A(inst_cellmath__61[12]), .B(inst_cellmath__61[13]));
NAND2XL inst_cellmath__203_0_I3993 (.Y(N12808), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
NOR2XL inst_cellmath__203_0_I3994 (.Y(N11882), .A(inst_cellmath__61[13]), .B(inst_cellmath__61[12]));
AND2XL inst_cellmath__203_0_I3995 (.Y(N13155), .A(N12808), .B(inst_cellmath__61[14]));
OR2XL inst_cellmath__203_0_I3996 (.Y(N11998), .A(N11882), .B(inst_cellmath__61[14]));
INVXL inst_cellmath__203_0_I3997 (.Y(N13225), .A(N13155));
NOR2XL inst_cellmath__203_0_I3998 (.Y(N12560), .A(N12763), .B(N12448));
MXI2XL inst_cellmath__203_0_I3999 (.Y(N12939), .A(N13225), .B(N11998), .S0(N12560));
MXI2XL inst_cellmath__203_0_I4000 (.Y(N12495), .A(N13123), .B(N12763), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4001 (.Y(N13324), .A(N13225), .B(N11998), .S0(N12495));
MXI2XL inst_cellmath__203_0_I4002 (.Y(N12430), .A(N11832), .B(N13123), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4003 (.Y(N12023), .A(N13225), .B(N11998), .S0(N12430));
MXI2XL inst_cellmath__203_0_I4004 (.Y(N12372), .A(N12203), .B(N11832), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4005 (.Y(N12384), .A(N13225), .B(N11998), .S0(N12372));
MXI2XL inst_cellmath__203_0_I4006 (.Y(N12310), .A(N12570), .B(N12203), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4007 (.Y(N12738), .A(N13225), .B(N11998), .S0(N12310));
MXI2XL inst_cellmath__203_0_I4008 (.Y(N12245), .A(N12905), .B(N12570), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4009 (.Y(N13093), .A(N13225), .B(N11998), .S0(N12245));
MXI2XL inst_cellmath__203_0_I4010 (.Y(N12185), .A(N13287), .B(N12905), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4011 (.Y(N11800), .A(N13225), .B(N11998), .S0(N12185));
MXI2XL inst_cellmath__203_0_I4012 (.Y(N12126), .A(N11992), .B(N13287), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4013 (.Y(N12171), .A(N13225), .B(N11998), .S0(N12126));
MXI2XL inst_cellmath__203_0_I4014 (.Y(N12065), .A(N12353), .B(N11992), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4015 (.Y(N12537), .A(N13225), .B(N11998), .S0(N12065));
MXI2XL inst_cellmath__203_0_I4016 (.Y(N12002), .A(N12708), .B(N12353), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4017 (.Y(N12874), .A(N13225), .B(N11998), .S0(N12002));
MXI2XL inst_cellmath__203_0_I4018 (.Y(N11936), .A(N13059), .B(N12708), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4019 (.Y(N13254), .A(N13225), .B(N11998), .S0(N11936));
MXI2XL inst_cellmath__203_0_I4020 (.Y(N11865), .A(N11770), .B(N13059), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4021 (.Y(N11963), .A(N13225), .B(N11998), .S0(N11865));
MXI2XL inst_cellmath__203_0_I4022 (.Y(N11804), .A(N12142), .B(N11770), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4023 (.Y(N12324), .A(N13225), .B(N11998), .S0(N11804));
MXI2XL inst_cellmath__203_0_I4024 (.Y(N11745), .A(N12507), .B(N12142), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4025 (.Y(N12684), .A(N13225), .B(N11998), .S0(N11745));
MXI2XL inst_cellmath__203_0_I4026 (.Y(N11680), .A(N12846), .B(N12507), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4027 (.Y(N13028), .A(N13225), .B(N11998), .S0(N11680));
MXI2XL inst_cellmath__203_0_I4028 (.Y(N13288), .A(N13218), .B(N12846), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4029 (.Y(N11738), .A(N13225), .B(N11998), .S0(N13288));
MXI2XL inst_cellmath__203_0_I4030 (.Y(N13219), .A(N11926), .B(N13218), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4031 (.Y(N12115), .A(N13225), .B(N11998), .S0(N13219));
MXI2XL inst_cellmath__203_0_I4032 (.Y(N13151), .A(N12292), .B(N11926), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4033 (.Y(N12477), .A(N13225), .B(N11998), .S0(N13151));
MXI2XL inst_cellmath__203_0_I4034 (.Y(N13088), .A(N12655), .B(N12292), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4035 (.Y(N12816), .A(N13225), .B(N11998), .S0(N13088));
MXI2XL inst_cellmath__203_0_I4036 (.Y(N13023), .A(N12996), .B(N12655), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4037 (.Y(N13186), .A(N13225), .B(N11998), .S0(N13023));
MXI2XL inst_cellmath__203_0_I4038 (.Y(N12962), .A(N11707), .B(N12996), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4039 (.Y(N11894), .A(N13225), .B(N11998), .S0(N12962));
MXI2XL inst_cellmath__203_0_I4040 (.Y(N12898), .A(N12084), .B(N11707), .S0(N12448));
MXI2XL inst_cellmath__203_0_I4041 (.Y(N12261), .A(N13225), .B(N11998), .S0(N12898));
NOR2BX1 inst_cellmath__203_0_I4042 (.Y(N12838), .AN(N12448), .B(N12084));
MXI2XL inst_cellmath__203_0_I4043 (.Y(N12719), .A(N13225), .B(N11998), .S0(N12838));
XNOR2X1 inst_cellmath__203_0_I4044 (.Y(N12412), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
NAND2XL inst_cellmath__203_0_I4045 (.Y(N12781), .A(inst_cellmath__61[15]), .B(inst_cellmath__61[14]));
NOR2XL inst_cellmath__203_0_I4046 (.Y(N11849), .A(inst_cellmath__61[14]), .B(inst_cellmath__61[15]));
AND2XL inst_cellmath__203_0_I4047 (.Y(N13121), .A(N12781), .B(inst_cellmath__115__W1[0]));
OR2XL inst_cellmath__203_0_I4048 (.Y(N12026), .A(N11849), .B(inst_cellmath__115__W1[0]));
INVXL inst_cellmath__203_0_I4049 (.Y(inst_cellmath__203__W0[42]), .A(N13121));
NOR2XL inst_cellmath__203_0_I4050 (.Y(N12528), .A(N12763), .B(N12412));
MXI2XL inst_cellmath__203_0_I4051 (.Y(N12903), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12528));
MXI2XL inst_cellmath__203_0_I4052 (.Y(N12465), .A(N13123), .B(N12763), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4053 (.Y(N13281), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12465));
MXI2XL inst_cellmath__203_0_I4054 (.Y(N12401), .A(N11832), .B(N13123), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4055 (.Y(N11987), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12401));
MXI2XL inst_cellmath__203_0_I4056 (.Y(N12340), .A(N12203), .B(N11832), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4057 (.Y(N12350), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12340));
MXI2XL inst_cellmath__203_0_I4058 (.Y(N12280), .A(N12570), .B(N12203), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4059 (.Y(N12704), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12280));
MXI2XL inst_cellmath__203_0_I4060 (.Y(N12218), .A(N12905), .B(N12570), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4061 (.Y(N13055), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12218));
MXI2XL inst_cellmath__203_0_I4062 (.Y(N12156), .A(N13287), .B(N12905), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4063 (.Y(N11766), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12156));
MXI2XL inst_cellmath__203_0_I4064 (.Y(N12097), .A(N11992), .B(N13287), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4065 (.Y(N12136), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12097));
MXI2XL inst_cellmath__203_0_I4066 (.Y(N12034), .A(N12353), .B(N11992), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4067 (.Y(N12503), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12034));
MXI2XL inst_cellmath__203_0_I4068 (.Y(N11972), .A(N12708), .B(N12353), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4069 (.Y(N12843), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N11972));
MXI2XL inst_cellmath__203_0_I4070 (.Y(N11902), .A(N13059), .B(N12708), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4071 (.Y(N13213), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N11902));
MXI2XL inst_cellmath__203_0_I4072 (.Y(N11837), .A(N11770), .B(N13059), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4073 (.Y(N11921), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N11837));
MXI2XL inst_cellmath__203_0_I4074 (.Y(N11776), .A(N12142), .B(N11770), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4075 (.Y(N12290), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N11776));
MXI2XL inst_cellmath__203_0_I4076 (.Y(N11712), .A(N12507), .B(N12142), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4077 (.Y(N12651), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N11712));
MXI2XL inst_cellmath__203_0_I4078 (.Y(N13325), .A(N12846), .B(N12507), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4079 (.Y(N12992), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N13325));
MXI2XL inst_cellmath__203_0_I4080 (.Y(N13257), .A(N13218), .B(N12846), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4081 (.Y(N11703), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N13257));
MXI2XL inst_cellmath__203_0_I4082 (.Y(N13188), .A(N11926), .B(N13218), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4083 (.Y(N12078), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N13188));
MXI2XL inst_cellmath__203_0_I4084 (.Y(N13122), .A(N12292), .B(N11926), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4085 (.Y(N12439), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N13122));
MXI2XL inst_cellmath__203_0_I4086 (.Y(N13057), .A(N12655), .B(N12292), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4087 (.Y(N12785), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N13057));
MXI2XL inst_cellmath__203_0_I4088 (.Y(N12994), .A(N12996), .B(N12655), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4089 (.Y(N13146), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12994));
MXI2XL inst_cellmath__203_0_I4090 (.Y(N12932), .A(N11707), .B(N12996), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4091 (.Y(N11854), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12932));
MXI2XL inst_cellmath__203_0_I4092 (.Y(N12869), .A(N12084), .B(N11707), .S0(N12412));
MXI2XL inst_cellmath__203_0_I4093 (.Y(N12225), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12869));
NOR2BX1 inst_cellmath__203_0_I4094 (.Y(N12810), .AN(N12412), .B(N12084));
MXI2XL inst_cellmath__203_0_I4095 (.Y(inst_cellmath__203__W1[42]), .A(inst_cellmath__203__W0[42]), .B(N12026), .S0(N12810));
ADDHX1 inst_cellmath__203_0_I4096 (.CO(N11845), .S(inst_cellmath__203__W0[1]), .A(inst_cellmath__198[19]), .B(N13299));
ADDHX1 inst_cellmath__203_0_I4097 (.CO(N12587), .S(inst_cellmath__203__W1[2]), .A(N12367), .B(N11845));
ADDHX1 inst_cellmath__203_0_I4098 (.CO(N13305), .S(N12924), .A(N13156), .B(N13069));
ADDFX1 inst_cellmath__203_0_I4099 (.CO(N12374), .S(inst_cellmath__203__W1[3]), .A(N12924), .B(N12766), .CI(N12587));
ADDFX1 inst_cellmath__203_0_I4100 (.CO(N13074), .S(inst_cellmath__203__W0[4]), .A(N12154), .B(N12602), .CI(N13128));
ADDFX1 inst_cellmath__203_0_I4101 (.CO(N12160), .S(inst_cellmath__203__W1[4]), .A(N13322), .B(N13305), .CI(N12374));
ADDFX1 inst_cellmath__203_0_I4102 (.CO(N12860), .S(N12523), .A(N13148), .B(N13327), .CI(inst_cellmath__61[2]));
ADDFX1 inst_cellmath__203_0_I4103 (.CO(N11941), .S(N13236), .A(N12856), .B(N12523), .CI(N12410));
ADDFX1 inst_cellmath__203_0_I4104 (.CO(N12670), .S(inst_cellmath__203__W0[5]), .A(N12024), .B(N11835), .CI(N12198));
ADDFX1 inst_cellmath__203_0_I4105 (.CO(inst_cellmath__203__W0[6]), .S(inst_cellmath__203__W1[5]), .A(N13074), .B(N13236), .CI(N12160));
ADDFX1 inst_cellmath__203_0_I4106 (.CO(N12460), .S(N12100), .A(N11857), .B(N12387), .CI(N12860));
ADDFX1 inst_cellmath__203_0_I4107 (.CO(N13169), .S(N12801), .A(N11939), .B(N12100), .CI(N12208));
ADDFX1 inst_cellmath__203_0_I4108 (.CO(N12247), .S(N11871), .A(N12568), .B(N11941), .CI(N12385));
ADDFXL inst_cellmath__203_0_I4109 (.CO(inst_cellmath__203__W0[7]), .S(inst_cellmath__203__W1[6]), .A(N12670), .B(N12801), .CI(N11871));
ADDFX1 inst_cellmath__203_0_I4110 (.CO(N12039), .S(N13332), .A(N13096), .B(N11671), .CI(N13116));
ADDFX1 inst_cellmath__203_0_I4111 (.CO(N12748), .S(N12396), .A(N13332), .B(N12227), .CI(N12460));
ADDFX1 inst_cellmath__203_0_I4112 (.CO(N11811), .S(N13106), .A(N12396), .B(N12665), .CI(N13312));
ADDFX1 inst_cellmath__203_0_I4113 (.CO(N12552), .S(N12187), .A(N12736), .B(N12574), .CI(N12901));
ADDFX1 inst_cellmath__203_0_I4114 (.CO(N13266), .S(N12886), .A(N13106), .B(N13083), .CI(N13169));
ADDFX1 inst_cellmath__203_0_I4115 (.CO(inst_cellmath__203__W0[8]), .S(inst_cellmath__203__W1[7]), .A(N12187), .B(N12247), .CI(N12886));
ADDFX1 inst_cellmath__203_0_I4116 (.CO(N13038), .S(N12694), .A(N11822), .B(N12175), .CI(N12595));
ADDFX1 inst_cellmath__203_0_I4117 (.CO(N12128), .S(N11749), .A(N12694), .B(N12039), .CI(N12748));
ADDFX1 inst_cellmath__203_0_I4118 (.CO(N12827), .S(N12488), .A(N11749), .B(N11719), .CI(N12908));
ADDFX1 inst_cellmath__203_0_I4119 (.CO(N11906), .S(N13197), .A(N13094), .B(N11811), .CI(N13282));
ADDFX1 inst_cellmath__203_0_I4120 (.CO(N12636), .S(N12273), .A(N12488), .B(N11792), .CI(N12552));
ADDFX1 inst_cellmath__203_0_I4121 (.CO(inst_cellmath__203__W0[9]), .S(inst_cellmath__203__W1[8]), .A(N13197), .B(N13266), .CI(N12273));
ADDFX1 inst_cellmath__203_0_I4122 (.CO(N12423), .S(N12067), .A(N12877), .B(N13307), .CI(N13077));
ADDFX1 inst_cellmath__203_0_I4123 (.CO(N13131), .S(N12773), .A(N12934), .B(N12195), .CI(N13038));
ADDFX1 inst_cellmath__203_0_I4124 (.CO(N12214), .S(N11840), .A(N12773), .B(N12067), .CI(N12454));
ADDFX1 inst_cellmath__203_0_I4125 (.CO(N12917), .S(N12578), .A(N12562), .B(N12128), .CI(N11840));
ADDFX1 inst_cellmath__203_0_I4126 (.CO(N12003), .S(N13296), .A(N12343), .B(N13291), .CI(N11801));
ADDFX1 inst_cellmath__203_0_I4127 (.CO(N12720), .S(N12364), .A(N12164), .B(N11988), .CI(N12578));
ADDFX1 inst_cellmath__203_0_I4128 (.CO(N11781), .S(N13066), .A(N11906), .B(N12827), .CI(N13296));
ADDFX1 inst_cellmath__203_0_I4129 (.CO(inst_cellmath__203__W0[10]), .S(inst_cellmath__203__W1[9]), .A(N12636), .B(N12364), .CI(N13066));
ADDFX1 inst_cellmath__203_0_I4130 (.CO(N13229), .S(N12854), .A(N11787), .B(N11965), .CI(N12564));
ADDFX1 inst_cellmath__203_0_I4131 (.CO(N12304), .S(N11937), .A(N12423), .B(N13316), .CI(N12854));
ADDFX1 inst_cellmath__203_0_I4132 (.CO(N13002), .S(N12664), .A(N11937), .B(N13131), .CI(N13161));
ADDFX1 inst_cellmath__203_0_I4133 (.CO(N12093), .S(N11716), .A(N12664), .B(N12214), .CI(N11997));
ADDFX1 inst_cellmath__203_0_I4134 (.CO(N12794), .S(N12451), .A(N12917), .B(N12700), .CI(N12172));
ADDFX1 inst_cellmath__203_0_I4135 (.CO(N11866), .S(N13160), .A(N12531), .B(N12348), .CI(N11716));
ADDFX1 inst_cellmath__203_0_I4136 (.CO(N12604), .S(N12236), .A(N12720), .B(N12003), .CI(N12451));
ADDFX1 inst_cellmath__203_0_I4137 (.CO(inst_cellmath__203__W0[11]), .S(inst_cellmath__203__W1[10]), .A(N11781), .B(N13160), .CI(N12236));
ADDFX1 inst_cellmath__203_0_I4138 (.CO(N12389), .S(N12030), .A(N12688), .B(N13268), .CI(N13040));
ADDFX1 inst_cellmath__203_0_I4139 (.CO(N13098), .S(N12741), .A(N12896), .B(N12162), .CI(N12016));
ADDFX1 inst_cellmath__203_0_I4140 (.CO(N12178), .S(N11805), .A(N12030), .B(N13229), .CI(N12741));
ADDFX1 inst_cellmath__203_0_I4141 (.CO(N12879), .S(N12544), .A(N12241), .B(N12304), .CI(N11805));
ADDFX1 inst_cellmath__203_0_I4142 (.CO(N11968), .S(N13259), .A(N11785), .B(N13002), .CI(N12544));
ADDFX1 inst_cellmath__203_0_I4143 (.CO(N12689), .S(N12328), .A(N13047), .B(N12356), .CI(N12538));
ADDFX1 inst_cellmath__203_0_I4144 (.CO(N11746), .S(N13032), .A(N12868), .B(N12705), .CI(N13233));
ADDFX1 inst_cellmath__203_0_I4145 (.CO(N12480), .S(N12120), .A(N13259), .B(N12093), .CI(N12794));
ADDFX1 inst_cellmath__203_0_I4146 (.CO(N13191), .S(N12820), .A(N13032), .B(N12328), .CI(N11866));
ADDFX1 inst_cellmath__203_0_I4147 (.CO(inst_cellmath__203__W0[12]), .S(inst_cellmath__203__W1[11]), .A(N12604), .B(N12120), .CI(N12820));
ADDFX1 inst_cellmath__203_0_I4148 (.CO(N12969), .S(N12629), .A(N11752), .B(N11743), .CI(N12526));
ADDFX1 inst_cellmath__203_0_I4149 (.CO(N12059), .S(N11681), .A(N12380), .B(N13277), .CI(N12389));
ADDFX1 inst_cellmath__203_0_I4150 (.CO(N12764), .S(N12416), .A(N12629), .B(N13098), .CI(N11681));
ADDFX1 inst_cellmath__203_0_I4151 (.CO(N11833), .S(N13124), .A(N12943), .B(N12178), .CI(N12416));
ADDFX1 inst_cellmath__203_0_I4152 (.CO(N12571), .S(N12204), .A(N12712), .B(N12879), .CI(N13124));
ADDFX1 inst_cellmath__203_0_I4153 (.CO(N13289), .S(N12907), .A(N12875), .B(N11757), .CI(N13056));
ADDFX1 inst_cellmath__203_0_I4154 (.CO(N12355), .S(N11993), .A(N11968), .B(N13243), .CI(N11942));
ADDFX1 inst_cellmath__203_0_I4155 (.CO(N13060), .S(N12709), .A(N12204), .B(N12689), .CI(N11746));
ADDFX1 inst_cellmath__203_0_I4156 (.CO(N12143), .S(N11771), .A(N11993), .B(N12907), .CI(N12480));
ADDFX1 inst_cellmath__203_0_I4157 (.CO(inst_cellmath__203__W0[13]), .S(inst_cellmath__203__W1[12]), .A(N13191), .B(N12709), .CI(N11771));
ADDFX1 inst_cellmath__203_0_I4158 (.CO(N11927), .S(N13220), .A(N12478), .B(N13230), .CI(N13004));
ADDFX1 inst_cellmath__203_0_I4159 (.CO(N12656), .S(N12295), .A(N12732), .B(N12130), .CI(N12862));
ADDFX1 inst_cellmath__203_0_I4160 (.CO(N11708), .S(N12997), .A(N12969), .B(N11983), .CI(N13220));
ADDFX1 inst_cellmath__203_0_I4161 (.CO(N12444), .S(N12087), .A(N12059), .B(N12295), .CI(N12997));
ADDFX1 inst_cellmath__203_0_I4162 (.CO(N13154), .S(N12789), .A(N12764), .B(N12032), .CI(N12087));
ADDFX1 inst_cellmath__203_0_I4163 (.CO(N12229), .S(N11859), .A(N12695), .B(N11833), .CI(N13063));
ADDFX1 inst_cellmath__203_0_I4164 (.CO(N12935), .S(N12599), .A(N12789), .B(N12133), .CI(N13255));
ADDFX1 inst_cellmath__203_0_I4165 (.CO(N12021), .S(N13319), .A(N11951), .B(N11764), .CI(N12311));
ADDFX1 inst_cellmath__203_0_I4166 (.CO(N12734), .S(N12381), .A(N12571), .B(N12487), .CI(N11859));
ADDFX1 inst_cellmath__203_0_I4167 (.CO(N11796), .S(N13092), .A(N12355), .B(N13289), .CI(N12599));
ADDFX1 inst_cellmath__203_0_I4168 (.CO(N12536), .S(N12169), .A(N13060), .B(N13319), .CI(N12381));
ADDFX1 inst_cellmath__203_0_I4169 (.CO(inst_cellmath__203__W0[14]), .S(inst_cellmath__203__W1[13]), .A(N13092), .B(N12143), .CI(N12169));
ADDFX1 inst_cellmath__203_0_I4170 (.CO(N12321), .S(N11959), .A(N11718), .B(N13190), .CI(N12491));
ADDFX1 inst_cellmath__203_0_I4171 (.CO(N13025), .S(N12682), .A(N13086), .B(N13238), .CI(N12344));
ADDFX1 inst_cellmath__203_0_I4172 (.CO(N12112), .S(N11735), .A(N12656), .B(N11927), .CI(N11959));
ADDFX1 inst_cellmath__203_0_I4173 (.CO(N12814), .S(N12474), .A(N11708), .B(N12682), .CI(N11735));
ADDFX1 inst_cellmath__203_0_I4174 (.CO(N11890), .S(N13183), .A(N12444), .B(N12746), .CI(N12474));
ADDFX1 inst_cellmath__203_0_I4175 (.CO(N12625), .S(N12259), .A(N13154), .B(N11773), .CI(N12496));
ADDFX1 inst_cellmath__203_0_I4176 (.CO(N11673), .S(N12964), .A(N12137), .B(N11961), .CI(N12317));
ADDFX1 inst_cellmath__203_0_I4177 (.CO(N12409), .S(N12051), .A(N12669), .B(N13183), .CI(N12828));
ADDFX1 inst_cellmath__203_0_I4178 (.CO(N13119), .S(N12759), .A(N12935), .B(N12229), .CI(N12021));
ADDFX1 inst_cellmath__203_0_I4179 (.CO(N12196), .S(N11826), .A(N12964), .B(N12259), .CI(N12734));
ADDFX1 inst_cellmath__203_0_I4180 (.CO(N12900), .S(N12566), .A(N11796), .B(N12051), .CI(N12759));
ADDFX1 inst_cellmath__203_0_I4181 (.CO(inst_cellmath__203__W0[15]), .S(inst_cellmath__203__W1[14]), .A(N12536), .B(N11826), .CI(N12566));
ADDHX1 inst_cellmath__203_0_I4182 (.CO(N12703), .S(N12347), .A(N13193), .B(N12265));
ADDFX1 inst_cellmath__203_0_I4183 (.CO(N11762), .S(N13052), .A(N12347), .B(N12971), .CI(N12096));
ADDFX1 inst_cellmath__203_0_I4184 (.CO(N12501), .S(N12135), .A(N12829), .B(N12702), .CI(N11944));
ADDFX1 inst_cellmath__203_0_I4185 (.CO(N13210), .S(N12840), .A(N12321), .B(N11794), .CI(N13025));
ADDFX1 inst_cellmath__203_0_I4186 (.CO(N12287), .S(N11918), .A(N12135), .B(N13052), .CI(N12112));
ADDFX1 inst_cellmath__203_0_I4187 (.CO(N12989), .S(N12649), .A(N11808), .B(N12840), .CI(N12814));
ADDFX1 inst_cellmath__203_0_I4188 (.CO(N12075), .S(N11699), .A(N13159), .B(N11918), .CI(N12146));
ADDFX1 inst_cellmath__203_0_I4189 (.CO(N12783), .S(N12437), .A(N12649), .B(N11890), .CI(N12833));
ADDFX1 inst_cellmath__203_0_I4190 (.CO(N11851), .S(N13143), .A(N12504), .B(N12325), .CI(N12676));
ADDFX1 inst_cellmath__203_0_I4191 (.CO(N12593), .S(N12223), .A(N13198), .B(N13008), .CI(N12625));
ADDFX1 inst_cellmath__203_0_I4192 (.CO(N13310), .S(N12930), .A(N11673), .B(N11699), .CI(N12437));
ADDFX1 inst_cellmath__203_0_I4193 (.CO(N12377), .S(N12011), .A(N13143), .B(N12409), .CI(N13119));
ADDFX1 inst_cellmath__203_0_I4194 (.CO(N13080), .S(N12729), .A(N12930), .B(N12223), .CI(N12196));
ADDFX1 inst_cellmath__203_0_I4195 (.CO(inst_cellmath__203__W0[16]), .S(inst_cellmath__203__W1[15]), .A(N12011), .B(N12900), .CI(N12729));
ADDFX1 inst_cellmath__203_0_I4196 (.CO(N12864), .S(N12529), .A(N12703), .B(N12966), .CI(N11684));
ADDFX1 inst_cellmath__203_0_I4197 (.CO(N11948), .S(N13241), .A(N13200), .B(N12453), .CI(N12313));
ADDFX1 inst_cellmath__203_0_I4198 (.CO(N12675), .S(N12314), .A(N12167), .B(N13050), .CI(N11762));
ADDFX1 inst_cellmath__203_0_I4199 (.CO(N11725), .S(N13015), .A(N12529), .B(N12501), .CI(N13241));
ADDFX1 inst_cellmath__203_0_I4200 (.CO(N12467), .S(N12103), .A(N12314), .B(N13210), .CI(N12545));
ADDFX1 inst_cellmath__203_0_I4201 (.CO(N13173), .S(N12805), .A(N12287), .B(N13015), .CI(N12103));
ADDFX1 inst_cellmath__203_0_I4202 (.CO(N12251), .S(N11880), .A(N12511), .B(N12989), .CI(N12237));
ADDFX1 inst_cellmath__203_0_I4203 (.CO(N12955), .S(N12617), .A(N12685), .B(N12841), .CI(N13205));
ADDFX1 inst_cellmath__203_0_I4204 (.CO(N12044), .S(N13337), .A(N12805), .B(N13017), .CI(N11722));
ADDFX1 inst_cellmath__203_0_I4205 (.CO(N12752), .S(N12404), .A(N12075), .B(N11904), .CI(N12783));
ADDFX1 inst_cellmath__203_0_I4206 (.CO(N11818), .S(N13109), .A(N11880), .B(N11851), .CI(N12617));
ADDFX1 inst_cellmath__203_0_I4207 (.CO(N12557), .S(N12190), .A(N12593), .B(N13337), .CI(N12404));
ADDFX1 inst_cellmath__203_0_I4208 (.CO(N13270), .S(N12891), .A(N13109), .B(N13310), .CI(N12377));
ADDFX1 inst_cellmath__203_0_I4209 (.CO(inst_cellmath__203__W0[17]), .S(inst_cellmath__203__W1[16]), .A(N13080), .B(N12190), .CI(N12891));
ADDFX1 inst_cellmath__203_0_I4210 (.CO(N13043), .S(N12698), .A(N12056), .B(N13155), .CI(N12939));
ADDFX1 inst_cellmath__203_0_I4211 (.CO(N12131), .S(N11756), .A(N12062), .B(N12533), .CI(N12673));
ADDFX1 inst_cellmath__203_0_I4212 (.CO(N12832), .S(N12493), .A(N11908), .B(N12797), .CI(N11760));
ADDFX1 inst_cellmath__203_0_I4213 (.CO(N11909), .S(N13202), .A(N12698), .B(N12864), .CI(N11948));
ADDFX1 inst_cellmath__203_0_I4214 (.CO(N12642), .S(N12281), .A(N12675), .B(N11756), .CI(N12493));
ADDFX1 inst_cellmath__203_0_I4215 (.CO(N11691), .S(N12981), .A(N13202), .B(N11725), .CI(N13263));
ADDFX1 inst_cellmath__203_0_I4216 (.CO(N12429), .S(N12070), .A(N12467), .B(N12281), .CI(N12981));
ADDFX1 inst_cellmath__203_0_I4217 (.CO(N13135), .S(N12776), .A(N12941), .B(N12848), .CI(N11912));
ADDFX1 inst_cellmath__203_0_I4218 (.CO(N12219), .S(N11843), .A(N13173), .B(N13026), .CI(N13214));
ADDFX1 inst_cellmath__203_0_I4219 (.CO(N12922), .S(N12585), .A(N12099), .B(N11729), .CI(N12070));
ADDFX1 inst_cellmath__203_0_I4220 (.CO(N12007), .S(N13302), .A(N12251), .B(N12274), .CI(N12955));
ADDFX1 inst_cellmath__203_0_I4221 (.CO(N12723), .S(N12371), .A(N12776), .B(N12044), .CI(N11843));
ADDFXL inst_cellmath__203_0_I4222 (.CO(N11783), .S(N13071), .A(N12585), .B(N12752), .CI(N13302));
ADDFX1 inst_cellmath__203_0_I4223 (.CO(N12520), .S(N12157), .A(N12371), .B(N11818), .CI(N12557));
ADDFX1 inst_cellmath__203_0_I4224 (.CO(inst_cellmath__203__W0[18]), .S(inst_cellmath__203__W1[17]), .A(N13270), .B(N13071), .CI(N12157));
ADDFX1 inst_cellmath__203_0_I4225 (.CO(N12308), .S(N11940), .A(N13324), .B(N12762), .CI(N12418));
ADDFX1 inst_cellmath__203_0_I4226 (.CO(N13006), .S(N12667), .A(N13163), .B(N12871), .CI(N12277));
ADDFX1 inst_cellmath__203_0_I4227 (.CO(N12098), .S(N11720), .A(N12134), .B(N13011), .CI(N13043));
ADDFX1 inst_cellmath__203_0_I4228 (.CO(N12799), .S(N12458), .A(N12832), .B(N12131), .CI(N11940));
ADDFX1 inst_cellmath__203_0_I4229 (.CO(N11870), .S(N13165), .A(N11720), .B(N12667), .CI(N11909));
ADDFXL inst_cellmath__203_0_I4230 (.CO(N12607), .S(N12243), .A(N12458), .B(N12332), .CI(N12642));
ADDFX1 inst_cellmath__203_0_I4231 (.CO(N13329), .S(N12946), .A(N11691), .B(N13165), .CI(N12243));
ADDFXL inst_cellmath__203_0_I4232 (.CO(N12394), .S(N12035), .A(N12029), .B(N13223), .CI(N12282));
ADDFX1 inst_cellmath__203_0_I4233 (.CO(N13102), .S(N12747), .A(N12429), .B(N11739), .CI(N11922));
ADDFX1 inst_cellmath__203_0_I4234 (.CO(N12183), .S(N11810), .A(N12461), .B(N12105), .CI(N12637));
ADDFXL inst_cellmath__203_0_I4235 (.CO(N12884), .S(N12549), .A(N12946), .B(N12219), .CI(N13135));
ADDFX1 inst_cellmath__203_0_I4236 (.CO(N11973), .S(N13264), .A(N12922), .B(N12035), .CI(N12747));
ADDFXL inst_cellmath__203_0_I4237 (.CO(N12693), .S(N12335), .A(N12007), .B(N11810), .CI(N12549));
ADDFX1 cynw_cm_float_cos_I29708 (.CO(N45668), .S(N13036), .A(N13264), .B(N12723), .CI(N11783));
ADDFX1 inst_cellmath__203_0_I4239 (.CO(inst_cellmath__203__W0[19]), .S(inst_cellmath__203__W1[18]), .A(N12520), .B(N12335), .CI(N13036));
ADDFX1 inst_cellmath__203_0_I4240 (.CO(N13195), .S(N12825), .A(N11830), .B(N13121), .CI(N12903));
ADDFX1 inst_cellmath__203_0_I4241 (.CO(N12271), .S(N11903), .A(N12023), .B(N12498), .CI(N12640));
ADDFX1 inst_cellmath__203_0_I4242 (.CO(N12973), .S(N12633), .A(N12765), .B(N13248), .CI(N11867));
ADDFX1 inst_cellmath__203_0_I4243 (.CO(N12064), .S(N11686), .A(N12308), .B(N11723), .CI(N12825));
ADDFX1 inst_cellmath__203_0_I4244 (.CO(N12770), .S(N12420), .A(N12098), .B(N13006), .CI(N11903));
ADDFX1 inst_cellmath__203_0_I4245 (.CO(N11839), .S(N13129), .A(N12799), .B(N12633), .CI(N11686));
ADDFX1 inst_cellmath__203_0_I4246 (.CO(N12575), .S(N12211), .A(N11870), .B(N13033), .CI(N12420));
ADDFXL inst_cellmath__203_0_I4247 (.CO(N13293), .S(N12913), .A(N13129), .B(N12607), .CI(N12211));
ADDFX1 inst_cellmath__203_0_I4248 (.CO(N12361), .S(N12000), .A(N11932), .B(N12742), .CI(N12644));
ADDFXL inst_cellmath__203_0_I4249 (.CO(N13064), .S(N12717), .A(N13329), .B(N12116), .CI(N12469));
ADDFX1 inst_cellmath__203_0_I4250 (.CO(N12150), .S(N11778), .A(N12975), .B(N12288), .CI(N12802));
ADDFXL inst_cellmath__203_0_I4251 (.CO(N12853), .S(N12512), .A(N12913), .B(N12394), .CI(N13102));
ADDFX1 inst_cellmath__203_0_I4252 (.CO(N11934), .S(N13227), .A(N12183), .B(N12000), .CI(N12717));
INVXL inst_cellmath__203_0_I4256 (.Y(N12757), .A(N12904));
ADDFX1 inst_cellmath__203_0_I4257 (.CO(N13158), .S(N12793), .A(N11954), .B(N12757), .CI(N13281));
ADDFX1 inst_cellmath__203_0_I4258 (.CO(N12940), .S(N12603), .A(N12384), .B(N13127), .CI(N12836));
ADDFX1 inst_cellmath__203_0_I4259 (.CO(N12027), .S(N13326), .A(N12240), .B(N12978), .CI(N12101));
ADDFX1 inst_cellmath__203_0_I4260 (.CO(N12740), .S(N12386), .A(N12271), .B(N13195), .CI(N12973));
ADDFX1 inst_cellmath__203_0_I4261 (.CO(N11803), .S(N13097), .A(N12793), .B(N12603), .CI(N13326));
ADDFX1 inst_cellmath__203_0_I4262 (.CO(N12541), .S(N12174), .A(N12770), .B(N12064), .CI(N12386));
ADDFX1 inst_cellmath__203_0_I4263 (.CO(N13258), .S(N12876), .A(N13097), .B(N23286), .CI(N11839));
ADDFX1 inst_cellmath__203_0_I4264 (.CO(N12326), .S(N11966), .A(N12174), .B(N12575), .CI(N12296));
ADDFX1 inst_cellmath__203_0_I4265 (.CO(N13029), .S(N12687), .A(N12876), .B(N11806), .CI(N12983));
ADDFXL inst_cellmath__203_0_I4266 (.CO(N12118), .S(N11742), .A(N12652), .B(N12475), .CI(N12809));
ADDFX1 inst_cellmath__203_0_I4267 (.CO(N12819), .S(N12479), .A(N13166), .B(N13293), .CI(N11687));
ADDFXL inst_cellmath__203_0_I4268 (.CO(N11896), .S(N13189), .A(N13064), .B(N11966), .CI(N12361));
ADDFX1 inst_cellmath__203_0_I4269 (.CO(N12628), .S(N12264), .A(N12150), .B(N12687), .CI(N11742));
ADDFX1 inst_cellmath__203_0_I4273 (.CO(N12202), .S(N11829), .A(N12319), .B(N13285), .CI(N12757));
ADDFX1 inst_cellmath__203_0_I4274 (.CO(N11990), .S(N13286), .A(N11987), .B(N12463), .CI(N12606));
ADDFX1 inst_cellmath__203_0_I4275 (.CO(N12707), .S(N12351), .A(N12738), .B(N13208), .CI(N11836));
ADDFX1 inst_cellmath__203_0_I4276 (.CO(N11768), .S(N13058), .A(N12940), .B(N11689), .CI(N13158));
ADDFX1 inst_cellmath__203_0_I4277 (.CO(N12505), .S(N12141), .A(N13286), .B(N12027), .CI(N11829));
ADDFX1 inst_cellmath__203_0_I4278 (.CO(N13217), .S(N12844), .A(N12740), .B(N12351), .CI(N13058));
ADDFXL inst_cellmath__203_0_I4279 (.CO(N12291), .S(N11924), .A(N12141), .B(N11803), .CI(N12541));
ADDFX1 inst_cellmath__203_0_I4280 (.CO(N12995), .S(N12654), .A(N13258), .B(N12844), .CI(N12659));
ADDFXL inst_cellmath__203_0_I4281 (.CO(N12083), .S(N11705), .A(N11924), .B(N12543), .CI(N11692));
ADDFX1 inst_cellmath__203_0_I4282 (.CO(N12786), .S(N12441), .A(N12817), .B(N12993), .CI(N13176));
ADDFX1 inst_cellmath__203_0_I4283 (.CO(N11856), .S(N13150), .A(N11872), .B(N12068), .CI(N12326));
ADDFXL inst_cellmath__203_0_I4284 (.CO(N12596), .S(N12226), .A(N12654), .B(N13029), .CI(N12118));
ADDFX1 inst_cellmath__203_0_I4285 (.CO(N13315), .S(N12933), .A(N12819), .B(N11705), .CI(N12441));
ADDFX1 inst_cellmath__203_0_I4289 (.CO(N12870), .S(N12534), .A(N12352), .B(N12904), .CI(N11916));
ADDFX1 inst_cellmath__203_0_I4290 (.CO(N11957), .S(N13247), .A(N13093), .B(N12350), .CI(N12804));
ADDFX1 inst_cellmath__203_0_I4291 (.CO(N12679), .S(N12318), .A(N12207), .B(N12942), .CI(N12069));
ADDFX1 inst_cellmath__203_0_I4292 (.CO(N11731), .S(N13022), .A(N11990), .B(N12680), .CI(N12202));
ADDFXL inst_cellmath__203_0_I4293 (.CO(N12472), .S(N12109), .A(N12534), .B(N12707), .CI(N13247));
ADDFX1 inst_cellmath__203_0_I4294 (.CO(N13180), .S(N12811), .A(N11768), .B(N12318), .CI(N13022));
ADDFX1 inst_cellmath__203_0_I4295 (.CO(N12256), .S(N11888), .A(N12109), .B(N12505), .CI(N13217));
ADDFX1 inst_cellmath__203_0_I4296 (.CO(N12961), .S(N12622), .A(N12725), .B(N12811), .CI(N12291));
ADDFXL inst_cellmath__203_0_I4297 (.CO(N12049), .S(N11670), .A(N13260), .B(N11888), .CI(N12071));
ADDFXL inst_cellmath__203_0_I4298 (.CO(N12758), .S(N12407), .A(N11701), .B(N13187), .CI(N11883));
ADDFX1 inst_cellmath__203_0_I4299 (.CO(N11824), .S(N13115), .A(N12424), .B(N12248), .CI(N12995));
ADDFXL inst_cellmath__203_0_I4300 (.CO(N12563), .S(N12194), .A(N12622), .B(N12083), .CI(N12786));
ADDFX1 inst_cellmath__203_0_I4301 (.CO(N13276), .S(N12897), .A(N12407), .B(N11670), .CI(N11856));
INVXL inst_cellmath__203_0_I4305 (.Y(N12646), .A(N11915));
ADDFX1 inst_cellmath__203_0_I4306 (.CO(N12837), .S(N12497), .A(N13170), .B(N12284), .CI(N12646));
ADDFX1 inst_cellmath__203_0_I4307 (.CO(N12647), .S(N12285), .A(N12573), .B(N12427), .CI(N12704));
ADDFX1 inst_cellmath__203_0_I4308 (.CO(N11696), .S(N12985), .A(N11800), .B(N13020), .CI(N13328));
ADDFX1 inst_cellmath__203_0_I4309 (.CO(N12433), .S(N12073), .A(N11957), .B(N12870), .CI(N12679));
ADDFX1 inst_cellmath__203_0_I4310 (.CO(N13142), .S(N12779), .A(N12497), .B(N12285), .CI(N12985));
ADDFXL inst_cellmath__203_0_I4311 (.CO(N12221), .S(N11848), .A(N12472), .B(N11731), .CI(N12073));
ADDFXL inst_cellmath__203_0_I4312 (.CO(N12927), .S(N12592), .A(N13180), .B(N12779), .CI(N11848));
ADDFXL inst_cellmath__203_0_I4313 (.CO(N12010), .S(N13306), .A(N12329), .B(N12256), .CI(N12432));
ADDFXL inst_cellmath__203_0_I4314 (.CO(N12727), .S(N12375), .A(N12079), .B(N11892), .CI(N12961));
ADDFXL inst_cellmath__203_0_I4315 (.CO(N11786), .S(N13078), .A(N12592), .B(N12255), .CI(N12610));
ADDFXL inst_cellmath__203_0_I4316 (.CO(N12527), .S(N12161), .A(N12771), .B(N12049), .CI(N12758));
ADDFXL inst_cellmath__203_0_I4317 (.CO(N13237), .S(N12861), .A(N12375), .B(N13306), .CI(N13078));
INVXL inst_cellmath__203_0_I4321 (.Y(N12589), .A(N11876));
ADDFX1 inst_cellmath__203_0_I4322 (.CO(N12803), .S(N12464), .A(N11875), .B(N11915), .CI(N12589));
ADDFX1 inst_cellmath__203_0_I4323 (.CO(N12613), .S(N12249), .A(N13055), .B(N12774), .CI(N12648));
ADDFX1 inst_cellmath__203_0_I4324 (.CO(N13334), .S(N12952), .A(N12910), .B(N11732), .CI(N12171));
ADDFX1 inst_cellmath__203_0_I4325 (.CO(N12400), .S(N12040), .A(N12837), .B(N12033), .CI(N12647));
ADDFX1 inst_cellmath__203_0_I4326 (.CO(N13107), .S(N12750), .A(N12464), .B(N11696), .CI(N12952));
ADDFX1 inst_cellmath__203_0_I4327 (.CO(N12189), .S(N11815), .A(N12433), .B(N12249), .CI(N12040));
ADDFX1 inst_cellmath__203_0_I4328 (.CO(N12889), .S(N12554), .A(N12750), .B(N13142), .CI(N12221));
ADDFXL inst_cellmath__203_0_I4329 (.CO(N11976), .S(N13267), .A(N12244), .B(N11815), .CI(N13031));
ADDFXL inst_cellmath__203_0_I4330 (.CO(N12696), .S(N12339), .A(N12927), .B(N12554), .CI(N12777));
ADDFX1 inst_cellmath__203_0_I4331 (.CO(N11753), .S(N13039), .A(N12619), .B(N12440), .CI(N12948));
ADDFXL inst_cellmath__203_0_I4332 (.CO(N12490), .S(N12129), .A(N13132), .B(N13267), .CI(N12010));
ADDFX1 inst_cellmath__203_0_I4333 (.CO(N13199), .S(N12830), .A(N11786), .B(N12727), .CI(N12339));
ADDFXL inst_cellmath__203_0_I4334 (.CO(N12279), .S(N11907), .A(N12527), .B(N13039), .CI(N12129));
ADDFXL cynw_cm_float_cos_I29584 (.CO(N12312), .S(N45350), .A(N11824), .B(N12563), .CI(N12161));
ADDFHXL inst_cellmath__203_0_I4335 (.CO(N12977), .S(N12639), .A(N12830), .B(N13237), .CI(N12312));
ADDFXL cynw_cm_float_cos_I29581 (.CO(N45345), .S(N45394), .A(N12596), .B(N13115), .CI(N12194));
ADDFXL cynw_cm_float_cos_I29585 (.CO(N13012), .S(N45377), .A(N12861), .B(N13276), .CI(N45345));
ADDFHXL inst_cellmath__203_0_I4336 (.CO(inst_cellmath__203__W0[25]), .S(inst_cellmath__203__W1[24]), .A(N13012), .B(N11907), .CI(N12639));
XNOR2X1 inst_cellmath__203_0_I4337 (.Y(N12426), .A(N12845), .B(N11876));
OR2XL inst_cellmath__203_0_I4338 (.Y(N12775), .A(N12845), .B(N11876));
ADDFX1 inst_cellmath__203_0_I4339 (.CO(N12582), .S(N12217), .A(N12250), .B(N12426), .CI(N12537));
ADDFX1 inst_cellmath__203_0_I4340 (.CO(N13300), .S(N12919), .A(N13133), .B(N12391), .CI(N12110));
ADDFX1 inst_cellmath__203_0_I4341 (.CO(N12368), .S(N12005), .A(N11766), .B(N12986), .CI(N13290));
ADDFX1 inst_cellmath__203_0_I4342 (.CO(N13068), .S(N12722), .A(N12613), .B(N12803), .CI(N13334));
ADDFX1 inst_cellmath__203_0_I4343 (.CO(N12155), .S(N11782), .A(N12919), .B(N12217), .CI(N12005));
ADDFX1 inst_cellmath__203_0_I4344 (.CO(N12857), .S(N12516), .A(N12400), .B(N13107), .CI(N12722));
ADDFX1 inst_cellmath__203_0_I4345 (.CO(N11938), .S(N13231), .A(N12189), .B(N11782), .CI(N12516));
ADDFXL inst_cellmath__203_0_I4346 (.CO(N12666), .S(N12306), .A(N12889), .B(N12121), .CI(N13138));
ADDFX1 inst_cellmath__203_0_I4347 (.CO(N11717), .S(N13003), .A(N12958), .B(N12784), .CI(N13333));
ADDFX1 inst_cellmath__203_0_I4348 (.CO(N12456), .S(N12095), .A(N11976), .B(N11841), .CI(N13231));
ADDFX1 inst_cellmath__203_0_I4349 (.CO(N13162), .S(N12796), .A(N11753), .B(N12696), .CI(N12306));
ADDFX1 inst_cellmath__203_0_I4350 (.CO(N12239), .S(N11869), .A(N12490), .B(N13003), .CI(N12095));
ADDFHXL inst_cellmath__203_0_I4351 (.CO(N12945), .S(N12605), .A(N12796), .B(N13199), .CI(N12279));
ADDFXL inst_cellmath__203_0_I4352 (.CO(inst_cellmath__203__W0[26]), .S(inst_cellmath__203__W1[25]), .A(N11869), .B(N12977), .CI(N12605));
ADDHX1 inst_cellmath__203_0_I4353 (.CO(N12744), .S(N12392), .A(N12775), .B(N12470));
ADDFX1 inst_cellmath__203_0_I4354 (.CO(N11809), .S(N13099), .A(N11842), .B(N12392), .CI(N12745));
ADDFX1 inst_cellmath__203_0_I4355 (.CO(N12546), .S(N12180), .A(N12874), .B(N11697), .CI(N12136));
ADDFX1 inst_cellmath__203_0_I4356 (.CO(N13261), .S(N12882), .A(N11996), .B(N12614), .CI(N12582));
ADDFX1 inst_cellmath__203_0_I4357 (.CO(N12333), .S(N11970), .A(N12368), .B(N13300), .CI(N13099));
ADDFX1 inst_cellmath__203_0_I4358 (.CO(N13034), .S(N12691), .A(N13068), .B(N12180), .CI(N12882));
ADDFX1 inst_cellmath__203_0_I4359 (.CO(N12123), .S(N11747), .A(N11970), .B(N12155), .CI(N12857));
ADDFX1 inst_cellmath__203_0_I4360 (.CO(N12823), .S(N12481), .A(N12125), .B(N12691), .CI(N12821));
ADDFX1 inst_cellmath__203_0_I4361 (.CO(N11901), .S(N13192), .A(N11938), .B(N11747), .CI(N11846));
ADDFXL inst_cellmath__203_0_I4362 (.CO(N12632), .S(N12269), .A(N12037), .B(N11668), .CI(N12213));
ADDFX1 inst_cellmath__203_0_I4363 (.CO(N11685), .S(N12970), .A(N12666), .B(N12481), .CI(N11717));
ADDFX1 inst_cellmath__203_0_I4364 (.CO(N12417), .S(N12061), .A(N12456), .B(N13192), .CI(N12269));
ADDFHXL inst_cellmath__203_0_I4365 (.CO(N13126), .S(N12768), .A(N12970), .B(N13162), .CI(N12239));
ADDFHXL inst_cellmath__203_0_I4366 (.CO(inst_cellmath__203__W0[27]), .S(inst_cellmath__203__W1[26]), .A(N12945), .B(N12061), .CI(N12768));
XNOR2X1 inst_cellmath__203_0_I4367 (.Y(N12572), .A(N12812), .B(N12744));
OR2XL inst_cellmath__203_0_I4368 (.Y(N12909), .A(N12812), .B(N12744));
ADDFX1 inst_cellmath__203_0_I4369 (.CO(N12714), .S(N12357), .A(N12216), .B(N12572), .CI(N12503));
ADDFX1 inst_cellmath__203_0_I4370 (.CO(N11774), .S(N13061), .A(N13100), .B(N12358), .CI(N12074));
ADDFX1 inst_cellmath__203_0_I4371 (.CO(N12509), .S(N12147), .A(N13254), .B(N12951), .CI(N11809));
ADDFX1 inst_cellmath__203_0_I4372 (.CO(N13224), .S(N12849), .A(N12357), .B(N12546), .CI(N13061));
ADDFX1 inst_cellmath__203_0_I4373 (.CO(N12297), .S(N11930), .A(N12333), .B(N13261), .CI(N12147));
ADDFX1 inst_cellmath__203_0_I4374 (.CO(N12999), .S(N12661), .A(N13034), .B(N12849), .CI(N11930));
ADDFX1 inst_cellmath__203_0_I4375 (.CO(N12088), .S(N11711), .A(N11898), .B(N12123), .CI(N12220));
ADDFXL inst_cellmath__203_0_I4376 (.CO(N12791), .S(N12447), .A(N12046), .B(N12661), .CI(N12397));
ADDFX1 inst_cellmath__203_0_I4377 (.CO(N11863), .S(N13157), .A(N12823), .B(N12579), .CI(N11901));
ADDFX1 inst_cellmath__203_0_I4378 (.CO(N12601), .S(N12232), .A(N12632), .B(N11711), .CI(N12447));
ADDFXL inst_cellmath__203_0_I4379 (.CO(N13323), .S(N12938), .A(N13157), .B(N11685), .CI(N12417));
ADDFXL inst_cellmath__203_0_I4380 (.CO(inst_cellmath__203__W0[28]), .S(inst_cellmath__203__W1[27]), .A(N13126), .B(N12232), .CI(N12938));
INVXL inst_cellmath__203_0_I4381 (.Y(N11874), .A(N10622));
ADDFX1 inst_cellmath__203_0_I4382 (.CO(N13095), .S(N12737), .A(N12434), .B(N11874), .CI(N12909));
ADDFX1 inst_cellmath__203_0_I4383 (.CO(N12873), .S(N12540), .A(N12711), .B(N11807), .CI(N13335));
ADDFX1 inst_cellmath__203_0_I4384 (.CO(N11962), .S(N13253), .A(N12583), .B(N12843), .CI(N11963));
ADDFX1 inst_cellmath__203_0_I4385 (.CO(N12683), .S(N12323), .A(N11774), .B(N12714), .CI(N12737));
ADDFX1 inst_cellmath__203_0_I4386 (.CO(N11740), .S(N13027), .A(N13253), .B(N12540), .CI(N12509));
ADDFX1 inst_cellmath__203_0_I4387 (.CO(N12476), .S(N12114), .A(N13224), .B(N12323), .CI(N13027));
ADDFX1 inst_cellmath__203_0_I4388 (.CO(N13185), .S(N12818), .A(N12297), .B(N12577), .CI(N12114));
ADDFX1 inst_cellmath__203_0_I4389 (.CO(N12263), .S(N11893), .A(N12630), .B(N12999), .CI(N12588));
ADDFX1 inst_cellmath__203_0_I4390 (.CO(N12965), .S(N12626), .A(N12918), .B(N12749), .CI(N12818));
ADDFX1 inst_cellmath__203_0_I4391 (.CO(N12053), .S(N11676), .A(N12791), .B(N12088), .CI(N11893));
ADDFXL inst_cellmath__203_0_I4392 (.CO(N12761), .S(N12411), .A(N12626), .B(N11863), .CI(N12601));
ADDFXL inst_cellmath__203_0_I4393 (.CO(inst_cellmath__203__W0[29]), .S(inst_cellmath__203__W1[28]), .A(N13323), .B(N11676), .CI(N12411));
ADDFX1 inst_cellmath__203_0_I4394 (.CO(N12567), .S(N12200), .A(N12181), .B(N12780), .CI(N10622));
ADDFX1 inst_cellmath__203_0_I4395 (.CO(N13283), .S(N12902), .A(N13062), .B(N12324), .CI(N12041));
ADDFXL inst_cellmath__203_0_I4396 (.CO(N12349), .S(N11986), .A(N13213), .B(N12920), .CI(N13095));
ADDFX1 inst_cellmath__203_0_I4397 (.CO(N13054), .S(N12706), .A(N12200), .B(N12873), .CI(N11962));
ADDFXL inst_cellmath__203_0_I4398 (.CO(N12139), .S(N11765), .A(N11986), .B(N12902), .CI(N12683));
ADDFXL inst_cellmath__203_0_I4399 (.CO(N12842), .S(N12502), .A(N11740), .B(N12706), .CI(N11765));
ADDFX1 inst_cellmath__203_0_I4400 (.CO(N11920), .S(N13215), .A(N12476), .B(N11682), .CI(N12502));
ADDFX1 inst_cellmath__203_0_I4401 (.CO(N12653), .S(N12289), .A(N13103), .B(N12925), .CI(N13185));
ADDFX1 inst_cellmath__203_0_I4402 (.CO(N11702), .S(N12991), .A(N12263), .B(N13295), .CI(N13215));
ADDFX1 inst_cellmath__203_0_I4403 (.CO(N12438), .S(N12081), .A(N12289), .B(N12965), .CI(N12053));
ADDFX1 inst_cellmath__203_0_I4404 (.CO(inst_cellmath__203__W0[30]), .S(inst_cellmath__203__W1[29]), .A(N12761), .B(N12991), .CI(N12081));
INVXL inst_cellmath__203_0_I4405 (.Y(N11814), .A(N12435));
ADDFX1 inst_cellmath__203_0_I4406 (.CO(N12224), .S(N11853), .A(N11775), .B(N12399), .CI(N11814));
ADDFX1 inst_cellmath__203_0_I4407 (.CO(N12015), .S(N13313), .A(N13298), .B(N12684), .CI(N12547));
ADDFX1 inst_cellmath__203_0_I4408 (.CO(N12730), .S(N12378), .A(N12567), .B(N11921), .CI(N13283));
ADDFX1 inst_cellmath__203_0_I4409 (.CO(N11791), .S(N13084), .A(N11853), .B(N12349), .CI(N13313));
ADDFX1 inst_cellmath__203_0_I4410 (.CO(N12532), .S(N12165), .A(N12378), .B(N13054), .CI(N12139));
ADDFX1 inst_cellmath__203_0_I4411 (.CO(N13244), .S(N12867), .A(N12165), .B(N13084), .CI(N11715));
ADDFX1 inst_cellmath__203_0_I4412 (.CO(N12316), .S(N11953), .A(N12415), .B(N12842), .CI(N11812));
ADDFX1 inst_cellmath__203_0_I4413 (.CO(N13018), .S(N12677), .A(N12867), .B(N12004), .CI(N11920));
ADDFXL inst_cellmath__203_0_I4414 (.CO(N12106), .S(N11728), .A(N11953), .B(N12653), .CI(N11702));
ADDFX1 inst_cellmath__203_0_I4415 (.CO(inst_cellmath__203__W0[31]), .S(inst_cellmath__203__W1[30]), .A(N12438), .B(N12677), .CI(N11728));
ADDFX1 inst_cellmath__203_0_I4416 (.CO(N11885), .S(N13177), .A(N12751), .B(N12435), .CI(N12145));
ADDFX1 inst_cellmath__203_0_I4417 (.CO(N12620), .S(N12254), .A(N13028), .B(N12290), .CI(N12006));
ADDFX1 inst_cellmath__203_0_I4418 (.CO(N11667), .S(N12959), .A(N12224), .B(N12880), .CI(N12015));
ADDFX1 inst_cellmath__203_0_I4419 (.CO(N12406), .S(N12047), .A(N12254), .B(N13177), .CI(N12730));
ADDFX1 inst_cellmath__203_0_I4420 (.CO(N13113), .S(N12756), .A(N12959), .B(N11791), .CI(N12047));
ADDFX1 inst_cellmath__203_0_I4421 (.CO(N12193), .S(N11821), .A(N12756), .B(N12532), .CI(N13125));
ADDFX1 inst_cellmath__203_0_I4422 (.CO(N12894), .S(N12561), .A(N12188), .B(N13244), .CI(N12365));
ADDFX1 inst_cellmath__203_0_I4423 (.CO(N11980), .S(N13275), .A(N12316), .B(N11821), .CI(N13018));
ADDFXL inst_cellmath__203_0_I4424 (.CO(inst_cellmath__203__W0[32]), .S(inst_cellmath__203__W1[31]), .A(N12106), .B(N12561), .CI(N13275));
INVXL inst_cellmath__203_0_I4425 (.Y(N11751), .A(N11877));
ADDFX1 inst_cellmath__203_0_I4426 (.CO(N11759), .S(N13046), .A(N11738), .B(N12369), .CI(N11751));
ADDFX1 inst_cellmath__203_0_I4427 (.CO(N13207), .S(N12834), .A(N13262), .B(N12651), .CI(N12510));
ADDFX1 inst_cellmath__203_0_I4428 (.CO(N12283), .S(N11911), .A(N12620), .B(N11885), .CI(N13046));
ADDFX1 inst_cellmath__203_0_I4429 (.CO(N12982), .S(N12645), .A(N11667), .B(N12834), .CI(N12406));
ADDFX1 inst_cellmath__203_0_I4430 (.CO(N12072), .S(N11694), .A(N13113), .B(N11911), .CI(N12645));
ADDFX1 inst_cellmath__203_0_I4431 (.CO(N12778), .S(N12431), .A(N12205), .B(N12177), .CI(N12718));
ADDFX1 inst_cellmath__203_0_I4432 (.CO(N11844), .S(N13140), .A(N12193), .B(N11694), .CI(N12894));
ADDFX1 inst_cellmath__203_0_I4433 (.CO(inst_cellmath__203__W0[33]), .S(inst_cellmath__203__W1[32]), .A(N11980), .B(N12431), .CI(N13140));
ADDFX1 inst_cellmath__203_0_I4434 (.CO(N13304), .S(N12923), .A(N12721), .B(N11877), .CI(N12115));
ADDFX1 inst_cellmath__203_0_I4435 (.CO(N12373), .S(N12008), .A(N11971), .B(N12992), .CI(N12850));
ADDFX1 inst_cellmath__203_0_I4436 (.CO(N13076), .S(N12726), .A(N13207), .B(N11759), .CI(N12923));
ADDFX1 inst_cellmath__203_0_I4437 (.CO(N12159), .S(N11784), .A(N12283), .B(N12008), .CI(N12726));
ADDFX1 inst_cellmath__203_0_I4438 (.CO(N12859), .S(N12524), .A(N11784), .B(N12982), .CI(N12906));
ADDFX1 inst_cellmath__203_0_I4439 (.CO(N11943), .S(N13235), .A(N13067), .B(N12072), .CI(N12524));
ADDFX1 inst_cellmath__203_0_I4440 (.CO(inst_cellmath__203__W1[34]), .S(inst_cellmath__203__W1[33]), .A(N11844), .B(N12778), .CI(N13235));
INVXL inst_cellmath__203_0_I4441 (.Y(N11688), .A(N12980));
ADDFX1 inst_cellmath__203_0_I4442 (.CO(N11721), .S(N13010), .A(N11703), .B(N12331), .CI(N11688));
ADDFX1 inst_cellmath__203_0_I4443 (.CO(N13168), .S(N12800), .A(N12477), .B(N13222), .CI(N13304));
ADDFX1 inst_cellmath__203_0_I4444 (.CO(N12246), .S(N11873), .A(N13010), .B(N12373), .CI(N12800));
ADDFX1 inst_cellmath__203_0_I4445 (.CO(N12950), .S(N12611), .A(N11873), .B(N13076), .CI(N12159));
ADDFX1 inst_cellmath__203_0_I4446 (.CO(N12038), .S(N13331), .A(N12611), .B(N11994), .CI(N12968));
ADDFX1 inst_cellmath__203_0_I4447 (.CO(inst_cellmath__203__W1[35]), .S(inst_cellmath__203__W0[34]), .A(N13331), .B(N12859), .CI(N11943));
ADDFX1 inst_cellmath__203_0_I4448 (.CO(N11813), .S(N13105), .A(N12692), .B(N12980), .CI(N12078));
ADDFX1 inst_cellmath__203_0_I4449 (.CO(N12551), .S(N12186), .A(N12816), .B(N11931), .CI(N11721));
ADDFX1 inst_cellmath__203_0_I4450 (.CO(N13265), .S(N12888), .A(N13168), .B(N13105), .CI(N12186));
ADDFX1 inst_cellmath__203_0_I4451 (.CO(N12337), .S(N11974), .A(N12888), .B(N12246), .CI(N12950));
ADDFX1 inst_cellmath__203_0_I4452 (.CO(inst_cellmath__203__W1[36]), .S(inst_cellmath__203__W0[35]), .A(N11974), .B(N12710), .CI(N12038));
INVXL inst_cellmath__203_0_I4453 (.Y(N13297), .A(N12457));
ADDFX1 inst_cellmath__203_0_I4454 (.CO(N12127), .S(N11750), .A(N13186), .B(N12298), .CI(N13297));
ADDFX1 inst_cellmath__203_0_I4455 (.CO(N11905), .S(N13196), .A(N11813), .B(N12439), .CI(N11750));
ADDFX1 inst_cellmath__203_0_I4456 (.CO(N12635), .S(N12275), .A(N13196), .B(N12551), .CI(N13265));
ADDFX1 inst_cellmath__203_0_I4457 (.CO(inst_cellmath__203__W1[37]), .S(inst_cellmath__203__W0[36]), .A(N13204), .B(N12275), .CI(N12337));
ADDFX1 inst_cellmath__203_0_I4458 (.CO(N12422), .S(N12066), .A(N12658), .B(N12457), .CI(N11894));
ADDFX1 inst_cellmath__203_0_I4459 (.CO(N13130), .S(N12772), .A(N12127), .B(N12785), .CI(N12066));
ADDFX1 inst_cellmath__203_0_I4460 (.CO(inst_cellmath__203__W1[38]), .S(inst_cellmath__203__W0[37]), .A(N12772), .B(N11905), .CI(N12635));
ADDFX1 inst_cellmath__203_0_I4461 (.CO(N12916), .S(N12581), .A(N12261), .B(N12484), .CI(N13146));
ADDFX1 inst_cellmath__203_0_I4462 (.CO(inst_cellmath__203__W1[39]), .S(inst_cellmath__203__W0[38]), .A(N12581), .B(N12422), .CI(N13130));
INVXL inst_cellmath__203_0_I4463 (.Y(N12363), .A(N12719));
ADDFX1 inst_cellmath__203_0_I4464 (.CO(inst_cellmath__203__W1[40]), .S(inst_cellmath__203__W0[39]), .A(N11854), .B(N12363), .CI(N12916));
ADDFX1 inst_cellmath__203_0_I4465 (.CO(inst_cellmath__203__W1[41]), .S(inst_cellmath__203__W0[40]), .A(N12719), .B(N13225), .CI(N12225));
INVXL inst_cellmath__203_0_I4466 (.Y(inst_cellmath__203__W0[41]), .A(inst_cellmath__203__W1[42]));
ADDHX1 cynw_cm_float_cos_I4469 (.CO(N15171), .S(N15033), .A(inst_cellmath__195[0]), .B(inst_cellmath__203__W0[18]));
ADDFXL cynw_cm_float_cos_I29709 (.CO(N45692), .S(N45679), .A(N12884), .B(N11778), .CI(N12512));
ADDFXL cynw_cm_float_cos_I29710 (.CO(N45718), .S(N45705), .A(N13227), .B(N11973), .CI(N12693));
ADDFXL cynw_cm_float_cos_I29711 (.CO(N45684), .S(inst_cellmath__203__W1[19]), .A(N45668), .B(N45679), .CI(N45705));
ADDFHX1 cynw_cm_float_cos_I4470 (.CO(N15461), .S(N15316), .A(inst_cellmath__195[1]), .B(inst_cellmath__203__W0[19]), .CI(inst_cellmath__203__W1[19]));
OR4X1 cynw_cm_float_cos_I30019 (.Y(N45720), .A(N8091), .B(N9030), .C(N9104), .D(N8038));
OR4X1 cynw_cm_float_cos_I30021 (.Y(N45700), .A(N8017), .B(N8290), .C(N8978), .D(N9056));
ADDFXL cynw_cm_float_cos_I29712 (.CO(N45711), .S(N45698), .A(N12479), .B(N12853), .CI(N13189));
ADDFXL cynw_cm_float_cos_I29713 (.CO(N45708), .S(N45695), .A(N12264), .B(N11934), .CI(N45692));
ADDFHXL cynw_cm_float_cos_I29714 (.CO(N45677), .S(N45724), .A(N45718), .B(N45698), .CI(N45695));
ADDFHX1 cynw_cm_float_cos_I29715 (.CO(N15089), .S(N14945), .A(N45720), .B(N45684), .CI(N45724));
ADDFXL cynw_cm_float_cos_I29716 (.CO(N45389), .S(N45721), .A(N11896), .B(N13150), .CI(N12226));
ADDFHXL cynw_cm_float_cos_I29717 (.CO(N45353), .S(N45687), .A(N12933), .B(N12628), .CI(N45711));
ADDFHXL cynw_cm_float_cos_I29718 (.CO(N45380), .S(N45713), .A(N45708), .B(N45721), .CI(N45687));
ADDFHX1 cynw_cm_float_cos_I29719 (.CO(N15373), .S(N15230), .A(N45677), .B(N45700), .CI(N45713));
NAND2X4 cynw_cm_float_cos_I29720 (.Y(N15196), .A(N15089), .B(N15230));
ADDFHXL cynw_cm_float_cos_I29582 (.CO(N45371), .S(N45358), .A(N13315), .B(N12897), .CI(N45389));
ADDFXL cynw_cm_float_cos_I29586 (.CO(inst_cellmath__203__W0[24]), .S(N45342), .A(N45371), .B(N45350), .CI(N45377));
ADDFHX1 cynw_cm_float_cos_I4475 (.CO(N15584), .S(N15433), .A(inst_cellmath__203__W0[24]), .B(inst_cellmath__195[6]), .CI(inst_cellmath__203__W1[24]));
ADDFHXL cynw_cm_float_cos_I4476 (.CO(N15205), .S(N15062), .A(inst_cellmath__195[7]), .B(inst_cellmath__203__W0[25]), .CI(inst_cellmath__203__W1[25]));
ADDFHXL cynw_cm_float_cos_I4477 (.CO(N15495), .S(N15349), .A(inst_cellmath__203__W0[26]), .B(inst_cellmath__195[8]), .CI(inst_cellmath__203__W1[26]));
ADDFX1 cynw_cm_float_cos_I4478 (.CO(N15124), .S(N14979), .A(inst_cellmath__203__W0[27]), .B(inst_cellmath__195[9]), .CI(inst_cellmath__203__W1[27]));
ADDFHXL cynw_cm_float_cos_I4479 (.CO(N15407), .S(N15262), .A(inst_cellmath__203__W0[28]), .B(inst_cellmath__195[10]), .CI(inst_cellmath__203__W1[28]));
ADDFHXL cynw_cm_float_cos_I4480 (.CO(N15041), .S(N15561), .A(inst_cellmath__203__W0[29]), .B(inst_cellmath__195[11]), .CI(inst_cellmath__203__W1[29]));
ADDFX1 cynw_cm_float_cos_I4481 (.CO(N15326), .S(N15182), .A(inst_cellmath__203__W0[30]), .B(inst_cellmath__195[12]), .CI(inst_cellmath__203__W1[30]));
ADDFX1 cynw_cm_float_cos_I4482 (.CO(N14954), .S(N15470), .A(inst_cellmath__203__W0[31]), .B(inst_cellmath__195[13]), .CI(inst_cellmath__203__W1[31]));
ADDFX1 cynw_cm_float_cos_I4483 (.CO(N15238), .S(N15101), .A(inst_cellmath__203__W0[32]), .B(inst_cellmath__195[14]), .CI(inst_cellmath__203__W1[32]));
ADDFX1 cynw_cm_float_cos_I4484 (.CO(N15535), .S(N15384), .A(inst_cellmath__203__W1[33]), .B(inst_cellmath__195[15]), .CI(inst_cellmath__203__W0[33]));
ADDFX1 cynw_cm_float_cos_I4485 (.CO(N15159), .S(N15016), .A(inst_cellmath__203__W0[34]), .B(inst_cellmath__195[16]), .CI(inst_cellmath__203__W1[34]));
ADDFX1 cynw_cm_float_cos_I4486 (.CO(N15445), .S(N15302), .A(inst_cellmath__203__W1[35]), .B(inst_cellmath__195[17]), .CI(inst_cellmath__203__W0[35]));
ADDFX1 cynw_cm_float_cos_I4487 (.CO(N15076), .S(N15595), .A(inst_cellmath__203__W0[36]), .B(inst_cellmath__195[18]), .CI(inst_cellmath__203__W1[36]));
ADDFX1 cynw_cm_float_cos_I4488 (.CO(N15359), .S(N15216), .A(inst_cellmath__203__W0[37]), .B(inst_cellmath__195[19]), .CI(inst_cellmath__203__W1[37]));
ADDFX1 cynw_cm_float_cos_I4489 (.CO(N14989), .S(N15509), .A(inst_cellmath__203__W0[38]), .B(inst_cellmath__195[20]), .CI(inst_cellmath__203__W1[38]));
ADDFX1 cynw_cm_float_cos_I4490 (.CO(N15274), .S(N15133), .A(inst_cellmath__203__W0[39]), .B(inst_cellmath__195[21]), .CI(inst_cellmath__203__W1[39]));
ADDFX1 cynw_cm_float_cos_I4491 (.CO(N15572), .S(N15417), .A(inst_cellmath__203__W0[40]), .B(inst_cellmath__195[22]), .CI(inst_cellmath__203__W1[40]));
ADDFX1 cynw_cm_float_cos_I4492 (.CO(N15191), .S(N15051), .A(inst_cellmath__195[23]), .B(inst_cellmath__203__W0[41]), .CI(inst_cellmath__203__W1[41]));
ADDFX1 cynw_cm_float_cos_I4493 (.CO(N15482), .S(N15335), .A(inst_cellmath__203__W1[42]), .B(inst_cellmath__203__W0[42]), .CI(inst_cellmath__195[24]));
ADDHX1 cynw_cm_float_cos_I4494 (.CO(N15111), .S(N14964), .A(1'B1), .B(inst_cellmath__195[25]));
ADDHX1 cynw_cm_float_cos_I4495 (.CO(N15394), .S(N15248), .A(1'B1), .B(inst_cellmath__195[26]));
ADDHX1 cynw_cm_float_cos_I4496 (.CO(N15027), .S(N15544), .A(1'B1), .B(inst_cellmath__195[27]));
INVXL hap1_A_I30022 (.Y(N15167), .A(inst_cellmath__195[28]));
OR2XL hap1_A_I11477 (.Y(N15313), .A(1'B0), .B(inst_cellmath__195[28]));
INVXL cynw_cm_float_cos_I4498 (.Y(N15455), .A(inst_cellmath__195[29]));
NOR2XL cynw_cm_float_cos_I4499 (.Y(N15519), .A(inst_cellmath__203__W0[1]), .B(inst_cellmath__203__W1[1]));
NOR2XL cynw_cm_float_cos_I4501 (.Y(N15144), .A(inst_cellmath__203__W0[2]), .B(inst_cellmath__203__W1[2]));
NAND2XL cynw_cm_float_cos_I4502 (.Y(N15284), .A(inst_cellmath__203__W0[2]), .B(inst_cellmath__203__W1[2]));
NOR2XL cynw_cm_float_cos_I4503 (.Y(N15429), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
NAND2XL cynw_cm_float_cos_I4504 (.Y(N15580), .A(inst_cellmath__203__W0[3]), .B(inst_cellmath__203__W1[3]));
AND2XL cynw_cm_float_cos_I4506 (.Y(N15201), .A(inst_cellmath__203__W0[4]), .B(inst_cellmath__203__W1[4]));
NOR2XL cynw_cm_float_cos_I4507 (.Y(N15345), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
NAND2XL cynw_cm_float_cos_I4508 (.Y(N15492), .A(inst_cellmath__203__W0[5]), .B(inst_cellmath__203__W1[5]));
NOR2XL cynw_cm_float_cos_I4509 (.Y(N14974), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
NAND2X1 cynw_cm_float_cos_I4510 (.Y(N15120), .A(inst_cellmath__203__W0[6]), .B(inst_cellmath__203__W1[6]));
OR2XL cynw_cm_float_cos_I4511 (.Y(N15257), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
AND2XL cynw_cm_float_cos_I4512 (.Y(N15403), .A(inst_cellmath__203__W0[7]), .B(inst_cellmath__203__W1[7]));
NOR2XL cynw_cm_float_cos_I4513 (.Y(N15556), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
NAND2XL cynw_cm_float_cos_I4514 (.Y(N15038), .A(inst_cellmath__203__W0[8]), .B(inst_cellmath__203__W1[8]));
OR2XL cynw_cm_float_cos_I4515 (.Y(N15177), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
AND2XL cynw_cm_float_cos_I4516 (.Y(N15322), .A(inst_cellmath__203__W0[9]), .B(inst_cellmath__203__W1[9]));
NOR2XL cynw_cm_float_cos_I4517 (.Y(N15466), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
NAND2XL cynw_cm_float_cos_I4518 (.Y(N14950), .A(inst_cellmath__203__W0[10]), .B(inst_cellmath__203__W1[10]));
NOR2XL cynw_cm_float_cos_I4519 (.Y(N15097), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
NAND2XL cynw_cm_float_cos_I4520 (.Y(N15234), .A(inst_cellmath__203__W0[11]), .B(inst_cellmath__203__W1[11]));
OR2XL cynw_cm_float_cos_I4521 (.Y(N15379), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
AND2XL cynw_cm_float_cos_I4522 (.Y(N15531), .A(inst_cellmath__203__W0[12]), .B(inst_cellmath__203__W1[12]));
NOR2XL cynw_cm_float_cos_I4523 (.Y(N15011), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NAND2XL cynw_cm_float_cos_I4524 (.Y(N15155), .A(inst_cellmath__203__W0[13]), .B(inst_cellmath__203__W1[13]));
NOR2XL cynw_cm_float_cos_I4525 (.Y(N15298), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NAND2XL cynw_cm_float_cos_I4526 (.Y(N15440), .A(inst_cellmath__203__W0[14]), .B(inst_cellmath__203__W1[14]));
NOR2XL cynw_cm_float_cos_I4527 (.Y(N15590), .A(inst_cellmath__203__W0[15]), .B(inst_cellmath__203__W1[15]));
NOR2XL cynw_cm_float_cos_I4529 (.Y(N15210), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
NAND2XL cynw_cm_float_cos_I4530 (.Y(N15355), .A(inst_cellmath__203__W0[16]), .B(inst_cellmath__203__W1[16]));
AOI21XL cynw_cm_float_cos_I4531 (.Y(N15129), .A0(N15284), .A1(N15519), .B0(N15144));
OAI2BB1X1 cynw_cm_float_cos_I10788 (.Y(N15270), .A0N(inst_cellmath__203__W0[1]), .A1N(inst_cellmath__203__W1[1]), .B0(N15284));
NAND2XL cynw_cm_float_cos_I4534 (.Y(N14960), .A(N15129), .B(N15270));
AOI21XL cynw_cm_float_cos_I4535 (.Y(N15453), .A0(N15580), .A1(N14960), .B0(N15429));
OAI22XL cynw_cm_float_cos_I10789 (.Y(N15199), .A0(N15201), .A1(N15453), .B0(inst_cellmath__203__W0[4]), .B1(inst_cellmath__203__W1[4]));
AO21XL cynw_cm_float_cos_I4539 (.Y(N14994), .A0(N15345), .A1(N15120), .B0(N14974));
AOI31X1 cynw_cm_float_cos_I4541 (.Y(N15068), .A0(N15120), .A1(N15492), .A2(N15199), .B0(N14994));
OAI21X1 cynw_cm_float_cos_I4544 (.Y(N15023), .A0(N15403), .A1(N15068), .B0(N15257));
AOI21X1 cynw_cm_float_cos_I4545 (.Y(N14970), .A0(N15038), .A1(N15023), .B0(N15556));
OAI21X1 cynw_cm_float_cos_I4548 (.Y(N15498), .A0(N15322), .A1(N14970), .B0(N15177));
AO21XL cynw_cm_float_cos_I4549 (.Y(N15327), .A0(N15466), .A1(N15234), .B0(N15097));
AOI31X2 cynw_cm_float_cos_I4551 (.Y(N15485), .A0(N15234), .A1(N14950), .A2(N15498), .B0(N15327));
OAI21X2 cynw_cm_float_cos_I4554 (.Y(N15560), .A0(N15531), .A1(N15485), .B0(N15379));
AO21XL cynw_cm_float_cos_I4555 (.Y(N15311), .A0(N15011), .A1(N15440), .B0(N15298));
AND2XL cynw_cm_float_cos_I4556 (.Y(N15456), .A(N15440), .B(N15155));
AOI21X2 cynw_cm_float_cos_I4560 (.Y(N15084), .A0(N15456), .A1(N15560), .B0(N15311));
AOI21XL cynw_cm_float_cos_I4563 (.Y(N15000), .A0(N15355), .A1(N15590), .B0(N15210));
OAI2BB1X1 cynw_cm_float_cos_I10794 (.Y(N15141), .A0N(inst_cellmath__203__W0[15]), .A1N(inst_cellmath__203__W1[15]), .B0(N15355));
OAI21X2 cynw_cm_float_cos_I4566 (.Y(N15598), .A0(N15141), .A1(N15084), .B0(N15000));
NOR2XL cynw_cm_float_cos_I4600 (.Y(N15221), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NAND2XL cynw_cm_float_cos_I4601 (.Y(N15362), .A(inst_cellmath__203__W0[17]), .B(inst_cellmath__203__W1[17]));
NOR2XL cynw_cm_float_cos_I4602 (.Y(N15514), .A(N15033), .B(inst_cellmath__203__W1[18]));
NAND2XL cynw_cm_float_cos_I4603 (.Y(N14995), .A(N15033), .B(inst_cellmath__203__W1[18]));
NOR2X2 cynw_cm_float_cos_I4604 (.Y(N15136), .A(N15171), .B(N15316));
NAND2X2 cynw_cm_float_cos_I4605 (.Y(N15279), .A(N15171), .B(N15316));
NOR2X2 cynw_cm_float_cos_I4606 (.Y(N15422), .A(N15461), .B(N14945));
NAND2X4 cynw_cm_float_cos_I4607 (.Y(N15574), .A(N15461), .B(N14945));
NOR2X2 cynw_cm_float_cos_I4608 (.Y(N15055), .A(N15089), .B(N15230));
OR4X1 cynw_cm_float_cos_I30030 (.Y(N45391), .A(N8976), .B(N8266), .C(N8263), .D(N8634));
ADDFHXL cynw_cm_float_cos_I29583 (.CO(N45400), .S(N45386), .A(N45353), .B(N45394), .CI(N45358));
ADDFHX1 cynw_cm_float_cos_I29587 (.CO(N15006), .S(N15522), .A(N45380), .B(N45391), .CI(N45386));
NOR2X2 cynw_cm_float_cos_I4610 (.Y(N15339), .A(N15373), .B(N15522));
NAND2X4 cynw_cm_float_cos_I4611 (.Y(N15488), .A(N15373), .B(N15522));
NOR2XL cynw_cm_float_cos_I29575 (.Y(N45383), .A(N8874), .B(N8758));
NOR2XL cynw_cm_float_cos_I29574 (.Y(N45368), .A(N9002), .B(N8084));
NOR2XL cynw_cm_float_cos_I29572 (.Y(N45341), .A(N8180), .B(N8824));
NOR2XL cynw_cm_float_cos_I29573 (.Y(N45355), .A(N9121), .B(N8159));
NAND4XL cynw_cm_float_cos_I29576 (.Y(N45397), .A(N45383), .B(N45368), .C(N45341), .D(N45355));
ADDFHX1 cynw_cm_float_cos_I29588 (.CO(N15288), .S(N15148), .A(N45400), .B(N45397), .CI(N45342));
NOR2X2 cynw_cm_float_cos_I4612 (.Y(N14968), .A(N15006), .B(N15148));
NAND2X4 cynw_cm_float_cos_I29589 (.Y(N15114), .A(N15006), .B(N15148));
NOR2X2 cynw_cm_float_cos_I4614 (.Y(N15254), .A(N15288), .B(N15433));
NAND2X4 cynw_cm_float_cos_I4615 (.Y(N15400), .A(N15288), .B(N15433));
NOR2X2 cynw_cm_float_cos_I4616 (.Y(N15549), .A(N15584), .B(N15062));
NAND2X2 cynw_cm_float_cos_I4617 (.Y(N15034), .A(N15584), .B(N15062));
NOR2X1 cynw_cm_float_cos_I4618 (.Y(N15173), .A(N15205), .B(N15349));
NAND2X2 cynw_cm_float_cos_I4619 (.Y(N15317), .A(N15205), .B(N15349));
NOR2X1 cynw_cm_float_cos_I4620 (.Y(N15462), .A(N15495), .B(N14979));
NAND2X2 cynw_cm_float_cos_I4621 (.Y(N14946), .A(N15495), .B(N14979));
NOR2X1 cynw_cm_float_cos_I4622 (.Y(N15090), .A(N15124), .B(N15262));
NAND2X2 cynw_cm_float_cos_I4623 (.Y(N15231), .A(N15124), .B(N15262));
NOR2X1 cynw_cm_float_cos_I4624 (.Y(N15374), .A(N15407), .B(N15561));
NAND2X1 cynw_cm_float_cos_I4625 (.Y(N15523), .A(N15561), .B(N15407));
NOR2X1 cynw_cm_float_cos_I4626 (.Y(N15007), .A(N15041), .B(N15182));
NAND2X2 cynw_cm_float_cos_I4627 (.Y(N15150), .A(N15041), .B(N15182));
NOR2XL cynw_cm_float_cos_I4628 (.Y(N15289), .A(N15326), .B(N15470));
NAND2X1 cynw_cm_float_cos_I4629 (.Y(N15434), .A(N15326), .B(N15470));
NOR2XL cynw_cm_float_cos_I4630 (.Y(N15585), .A(N14954), .B(N15101));
NAND2X1 cynw_cm_float_cos_I4631 (.Y(N15063), .A(N14954), .B(N15101));
NOR2XL cynw_cm_float_cos_I4632 (.Y(N15206), .A(N15384), .B(N15238));
NAND2XL cynw_cm_float_cos_I4633 (.Y(N15350), .A(N15384), .B(N15238));
NOR2XL cynw_cm_float_cos_I4634 (.Y(N15496), .A(N15535), .B(N15016));
NAND2XL cynw_cm_float_cos_I4635 (.Y(N14980), .A(N15535), .B(N15016));
NOR2XL cynw_cm_float_cos_I4636 (.Y(N15125), .A(N15159), .B(N15302));
NAND2XL cynw_cm_float_cos_I4637 (.Y(N15263), .A(N15159), .B(N15302));
NOR2XL cynw_cm_float_cos_I4638 (.Y(N15408), .A(N15595), .B(N15445));
NAND2XL cynw_cm_float_cos_I4639 (.Y(N15563), .A(N15595), .B(N15445));
NOR2XL cynw_cm_float_cos_I4640 (.Y(N15042), .A(N15216), .B(N15076));
NAND2XL cynw_cm_float_cos_I4641 (.Y(N15183), .A(N15216), .B(N15076));
NOR2XL cynw_cm_float_cos_I4642 (.Y(N15328), .A(N15509), .B(N15359));
NAND2XL cynw_cm_float_cos_I4643 (.Y(N15471), .A(N15509), .B(N15359));
NOR2XL cynw_cm_float_cos_I4644 (.Y(N14955), .A(N15133), .B(N14989));
NAND2XL cynw_cm_float_cos_I4645 (.Y(N15103), .A(N15133), .B(N14989));
NOR2XL cynw_cm_float_cos_I4646 (.Y(N15239), .A(N15417), .B(N15274));
NAND2XL cynw_cm_float_cos_I4647 (.Y(N15385), .A(N15417), .B(N15274));
NOR2XL cynw_cm_float_cos_I4648 (.Y(N15536), .A(N15051), .B(N15572));
NAND2XL cynw_cm_float_cos_I4649 (.Y(N15017), .A(N15051), .B(N15572));
NOR2XL cynw_cm_float_cos_I4650 (.Y(N15160), .A(N15335), .B(N15191));
NAND2XL cynw_cm_float_cos_I4651 (.Y(N15304), .A(N15335), .B(N15191));
NOR2XL cynw_cm_float_cos_I4652 (.Y(N15446), .A(N15482), .B(N14964));
NAND2XL cynw_cm_float_cos_I4653 (.Y(N15596), .A(N15482), .B(N14964));
NOR2XL cynw_cm_float_cos_I4654 (.Y(N15079), .A(N15111), .B(N15248));
NAND2XL cynw_cm_float_cos_I4655 (.Y(N15217), .A(N15111), .B(N15248));
NOR2XL cynw_cm_float_cos_I4656 (.Y(N15360), .A(N15544), .B(N15394));
NAND2XL cynw_cm_float_cos_I4657 (.Y(N15511), .A(N15544), .B(N15394));
NOR2XL cynw_cm_float_cos_I4658 (.Y(N14990), .A(N15167), .B(N15027));
NAND2XL cynw_cm_float_cos_I4659 (.Y(N15134), .A(N15167), .B(N15027));
NOR2XL cynw_cm_float_cos_I4660 (.Y(N15276), .A(N15455), .B(N15313));
NAND2XL cynw_cm_float_cos_I4661 (.Y(N15418), .A(N15455), .B(N15313));
INVXL cynw_cm_float_cos_I4662 (.Y(N14949), .A(N15598));
AOI21X1 cynw_cm_float_cos_I4663 (.Y(N15336), .A0(N15362), .A1(N15598), .B0(N15221));
AOI21X1 cynw_cm_float_cos_I4664 (.Y(N14965), .A0(N14995), .A1(N15221), .B0(N15514));
NAND2XL cynw_cm_float_cos_I4665 (.Y(N15112), .A(N14995), .B(N15362));
AOI21X2 cynw_cm_float_cos_I4666 (.Y(N15250), .A0(N15279), .A1(N15514), .B0(N15136));
NAND2XL cynw_cm_float_cos_I4667 (.Y(N15395), .A(N14995), .B(N15279));
AOI21X4 cynw_cm_float_cos_I4668 (.Y(N15546), .A0(N15136), .A1(N15574), .B0(N15422));
NAND2X2 cynw_cm_float_cos_I4669 (.Y(N15029), .A(N15279), .B(N15574));
AOI21X4 cynw_cm_float_cos_I4670 (.Y(N15168), .A0(N15196), .A1(N15422), .B0(N15055));
NAND2X2 cynw_cm_float_cos_I4671 (.Y(N15315), .A(N15196), .B(N15574));
AOI21X4 cynw_cm_float_cos_I4672 (.Y(N15458), .A0(N15488), .A1(N15055), .B0(N15339));
NAND2X2 cynw_cm_float_cos_I4673 (.Y(N14942), .A(N15488), .B(N15196));
AOI21X2 cynw_cm_float_cos_I4674 (.Y(N15088), .A0(N15114), .A1(N15339), .B0(N14968));
NAND2X2 cynw_cm_float_cos_I4675 (.Y(N15227), .A(N15488), .B(N15114));
AOI21X4 cynw_cm_float_cos_I4676 (.Y(N15370), .A0(N14968), .A1(N15400), .B0(N15254));
NAND2X4 cynw_cm_float_cos_I4677 (.Y(N15521), .A(N15400), .B(N15114));
AOI21X2 cynw_cm_float_cos_I4678 (.Y(N15003), .A0(N15034), .A1(N15254), .B0(N15549));
NAND2X2 cynw_cm_float_cos_I4679 (.Y(N15145), .A(N15034), .B(N15400));
AOI21X4 cynw_cm_float_cos_I4680 (.Y(N15286), .A0(N15317), .A1(N15549), .B0(N15173));
NAND2X2 cynw_cm_float_cos_I4681 (.Y(N15430), .A(N15317), .B(N15034));
AOI21X2 cynw_cm_float_cos_I4682 (.Y(N15581), .A0(N15173), .A1(N14946), .B0(N15462));
NAND2X2 cynw_cm_float_cos_I4683 (.Y(N15061), .A(N14946), .B(N15317));
AOI21X2 cynw_cm_float_cos_I4684 (.Y(N15202), .A0(N15231), .A1(N15462), .B0(N15090));
NAND2X2 cynw_cm_float_cos_I4685 (.Y(N15346), .A(N15231), .B(N14946));
AOI21X1 cynw_cm_float_cos_I4686 (.Y(N15494), .A0(N15523), .A1(N15090), .B0(N15374));
NAND2X1 cynw_cm_float_cos_I4687 (.Y(N14975), .A(N15231), .B(N15523));
AOI21X1 cynw_cm_float_cos_I4688 (.Y(N15121), .A0(N15374), .A1(N15150), .B0(N15007));
NAND2X1 cynw_cm_float_cos_I4689 (.Y(N15260), .A(N15150), .B(N15523));
AOI21X1 cynw_cm_float_cos_I4690 (.Y(N15404), .A0(N15434), .A1(N15007), .B0(N15289));
NAND2X1 cynw_cm_float_cos_I4691 (.Y(N15557), .A(N15434), .B(N15150));
AOI21XL cynw_cm_float_cos_I4692 (.Y(N15039), .A0(N15063), .A1(N15289), .B0(N15585));
NAND2X1 cynw_cm_float_cos_I4693 (.Y(N15178), .A(N15063), .B(N15434));
AOI21XL cynw_cm_float_cos_I4694 (.Y(N15323), .A0(N15350), .A1(N15585), .B0(N15206));
NAND2XL cynw_cm_float_cos_I4695 (.Y(N15467), .A(N15350), .B(N15063));
AOI21XL cynw_cm_float_cos_I4696 (.Y(N14951), .A0(N14980), .A1(N15206), .B0(N15496));
NAND2XL cynw_cm_float_cos_I4697 (.Y(N15099), .A(N14980), .B(N15350));
AOI21XL cynw_cm_float_cos_I4698 (.Y(N15236), .A0(N15263), .A1(N15496), .B0(N15125));
NAND2XL cynw_cm_float_cos_I4699 (.Y(N15380), .A(N15263), .B(N14980));
AOI21XL cynw_cm_float_cos_I4700 (.Y(N15533), .A0(N15563), .A1(N15125), .B0(N15408));
NAND2XL cynw_cm_float_cos_I4701 (.Y(N15013), .A(N15563), .B(N15263));
AOI21XL cynw_cm_float_cos_I4702 (.Y(N15156), .A0(N15183), .A1(N15408), .B0(N15042));
NAND2XL cynw_cm_float_cos_I4703 (.Y(N15300), .A(N15183), .B(N15563));
AOI21XL cynw_cm_float_cos_I4704 (.Y(N15442), .A0(N15471), .A1(N15042), .B0(N15328));
NAND2XL cynw_cm_float_cos_I4705 (.Y(N15591), .A(N15471), .B(N15183));
AOI21XL cynw_cm_float_cos_I4706 (.Y(N15074), .A0(N15103), .A1(N15328), .B0(N14955));
NAND2XL cynw_cm_float_cos_I4707 (.Y(N15212), .A(N15103), .B(N15471));
AOI21XL cynw_cm_float_cos_I4708 (.Y(N15356), .A0(N15385), .A1(N14955), .B0(N15239));
NAND2XL cynw_cm_float_cos_I4709 (.Y(N15507), .A(N15385), .B(N15103));
AOI21XL cynw_cm_float_cos_I4710 (.Y(N14986), .A0(N15017), .A1(N15239), .B0(N15536));
NAND2XL cynw_cm_float_cos_I4711 (.Y(N15130), .A(N15017), .B(N15385));
AOI21XL cynw_cm_float_cos_I4712 (.Y(N15272), .A0(N15304), .A1(N15536), .B0(N15160));
NAND2XL cynw_cm_float_cos_I4713 (.Y(N15413), .A(N15304), .B(N15017));
AOI21XL cynw_cm_float_cos_I4714 (.Y(N15568), .A0(N15596), .A1(N15160), .B0(N15446));
NAND2XL cynw_cm_float_cos_I4715 (.Y(N15049), .A(N15596), .B(N15304));
AOI21XL cynw_cm_float_cos_I4716 (.Y(N15188), .A0(N15217), .A1(N15446), .B0(N15079));
NAND2XL cynw_cm_float_cos_I4717 (.Y(N15332), .A(N15217), .B(N15596));
AOI21XL cynw_cm_float_cos_I4718 (.Y(N15480), .A0(N15511), .A1(N15079), .B0(N15360));
NAND2XL cynw_cm_float_cos_I4719 (.Y(N14961), .A(N15511), .B(N15217));
AOI21XL cynw_cm_float_cos_I4720 (.Y(N15108), .A0(N15134), .A1(N15360), .B0(N14990));
NAND2XL cynw_cm_float_cos_I4721 (.Y(N15246), .A(N15134), .B(N15511));
AOI21XL cynw_cm_float_cos_I4722 (.Y(N15391), .A0(N15418), .A1(N14990), .B0(N15276));
NAND2XL cynw_cm_float_cos_I4723 (.Y(N15541), .A(N15418), .B(N15134));
NAND2XL cynw_cm_float_cos_I4724 (.Y(N15309), .A(N15455), .B(N15418));
INVXL cynw_cm_float_cos_I4725 (.Y(N15096), .A(N14949));
INVXL cynw_cm_float_cos_I4726 (.Y(N15235), .A(N15336));
OAI21X1 cynw_cm_float_cos_I4727 (.Y(N15367), .A0(N15112), .A1(N14949), .B0(N14965));
OAI21X1 cynw_cm_float_cos_I4728 (.Y(N14999), .A0(N15395), .A1(N15336), .B0(N15250));
OAI21X2 cynw_cm_float_cos_I4729 (.Y(N15281), .A0(N14965), .A1(N15029), .B0(N15546));
NOR2X2 cynw_cm_float_cos_I4730 (.Y(N15427), .A(N15112), .B(N15029));
OAI21X2 cynw_cm_float_cos_I4731 (.Y(N15578), .A0(N15315), .A1(N15250), .B0(N15168));
NOR2X1 cynw_cm_float_cos_I4732 (.Y(N15057), .A(N15315), .B(N15395));
OAI21X1 cynw_cm_float_cos_I4733 (.Y(N15200), .A0(N14942), .A1(N15546), .B0(N15458));
NOR2X1 cynw_cm_float_cos_I4734 (.Y(N15343), .A(N15029), .B(N14942));
OAI21X2 cynw_cm_float_cos_I4735 (.Y(N15490), .A0(N15227), .A1(N15168), .B0(N15088));
NOR2X1 cynw_cm_float_cos_I4736 (.Y(N14973), .A(N15315), .B(N15227));
OAI21X4 cynw_cm_float_cos_I4737 (.Y(N15117), .A0(N15521), .A1(N15458), .B0(N15370));
NOR2X2 cynw_cm_float_cos_I4738 (.Y(N15255), .A(N14942), .B(N15521));
OAI21X2 cynw_cm_float_cos_I4739 (.Y(N15402), .A0(N15145), .A1(N15088), .B0(N15003));
NOR2X1 cynw_cm_float_cos_I4740 (.Y(N15554), .A(N15227), .B(N15145));
OAI21X2 cynw_cm_float_cos_I4741 (.Y(N15036), .A0(N15430), .A1(N15370), .B0(N15286));
NOR2X1 cynw_cm_float_cos_I4742 (.Y(N15176), .A(N15430), .B(N15521));
OAI21X2 cynw_cm_float_cos_I4743 (.Y(N15320), .A0(N15061), .A1(N15003), .B0(N15581));
NOR2X1 cynw_cm_float_cos_I4744 (.Y(N15464), .A(N15061), .B(N15145));
OAI21X4 cynw_cm_float_cos_I4745 (.Y(N14948), .A0(N15346), .A1(N15286), .B0(N15202));
NOR2X4 cynw_cm_float_cos_I4746 (.Y(N15094), .A(N15346), .B(N15430));
OAI21X2 cynw_cm_float_cos_I4747 (.Y(N15232), .A0(N14975), .A1(N15581), .B0(N15494));
NOR2X1 cynw_cm_float_cos_I4748 (.Y(N15377), .A(N14975), .B(N15061));
OAI21X1 cynw_cm_float_cos_I4749 (.Y(N15528), .A0(N15260), .A1(N15202), .B0(N15121));
NOR2X1 cynw_cm_float_cos_I4750 (.Y(N15009), .A(N15260), .B(N15346));
OAI21X1 cynw_cm_float_cos_I4751 (.Y(N15153), .A0(N15557), .A1(N15494), .B0(N15404));
NOR2X1 cynw_cm_float_cos_I4752 (.Y(N15295), .A(N15557), .B(N14975));
OAI21X1 cynw_cm_float_cos_I4753 (.Y(N15437), .A0(N15178), .A1(N15121), .B0(N15039));
NOR2X2 cynw_cm_float_cos_I4754 (.Y(N15588), .A(N15178), .B(N15260));
OAI21X1 cynw_cm_float_cos_I4755 (.Y(N15069), .A0(N15467), .A1(N15404), .B0(N15323));
NOR2X1 cynw_cm_float_cos_I4756 (.Y(N15208), .A(N15467), .B(N15557));
OAI21X1 cynw_cm_float_cos_I4757 (.Y(N15353), .A0(N15099), .A1(N15039), .B0(N14951));
NOR2X1 cynw_cm_float_cos_I4758 (.Y(N15503), .A(N15099), .B(N15178));
OAI21XL cynw_cm_float_cos_I4759 (.Y(N14982), .A0(N15380), .A1(N15323), .B0(N15236));
NOR2XL cynw_cm_float_cos_I4760 (.Y(N15128), .A(N15380), .B(N15467));
OAI21XL cynw_cm_float_cos_I4761 (.Y(N15268), .A0(N15013), .A1(N14951), .B0(N15533));
NOR2XL cynw_cm_float_cos_I4762 (.Y(N15410), .A(N15013), .B(N15099));
OAI21XL cynw_cm_float_cos_I4763 (.Y(N15566), .A0(N15300), .A1(N15236), .B0(N15156));
NOR2XL cynw_cm_float_cos_I4764 (.Y(N15047), .A(N15300), .B(N15380));
OAI21XL cynw_cm_float_cos_I4765 (.Y(N15185), .A0(N15591), .A1(N15533), .B0(N15442));
NOR2XL cynw_cm_float_cos_I4766 (.Y(N15331), .A(N15591), .B(N15013));
OAI21XL cynw_cm_float_cos_I4767 (.Y(N15477), .A0(N15212), .A1(N15156), .B0(N15074));
NOR2XL cynw_cm_float_cos_I4768 (.Y(N14957), .A(N15212), .B(N15300));
OAI21XL cynw_cm_float_cos_I4769 (.Y(N15106), .A0(N15507), .A1(N15442), .B0(N15356));
NOR2XL cynw_cm_float_cos_I4770 (.Y(N15244), .A(N15507), .B(N15591));
OAI21XL cynw_cm_float_cos_I4771 (.Y(N15387), .A0(N15130), .A1(N15074), .B0(N14986));
NOR2XL cynw_cm_float_cos_I4772 (.Y(N15540), .A(N15130), .B(N15212));
OAI21XL cynw_cm_float_cos_I4773 (.Y(N15024), .A0(N15413), .A1(N15356), .B0(N15272));
NOR2XL cynw_cm_float_cos_I4774 (.Y(N15162), .A(N15413), .B(N15507));
OAI21XL cynw_cm_float_cos_I4775 (.Y(N15307), .A0(N15049), .A1(N14986), .B0(N15568));
NOR2XL cynw_cm_float_cos_I4776 (.Y(N15451), .A(N15049), .B(N15130));
OAI21XL cynw_cm_float_cos_I4777 (.Y(N15599), .A0(N15332), .A1(N15272), .B0(N15188));
NOR2XL cynw_cm_float_cos_I4778 (.Y(N15082), .A(N15332), .B(N15413));
OAI21XL cynw_cm_float_cos_I4779 (.Y(N15223), .A0(N14961), .A1(N15568), .B0(N15480));
NOR2XL cynw_cm_float_cos_I4780 (.Y(N15363), .A(N14961), .B(N15049));
OAI21XL cynw_cm_float_cos_I4781 (.Y(N15515), .A0(N15246), .A1(N15188), .B0(N15108));
NOR2XL cynw_cm_float_cos_I4782 (.Y(N14997), .A(N15246), .B(N15332));
OAI21XL cynw_cm_float_cos_I4783 (.Y(N15137), .A0(N15541), .A1(N15480), .B0(N15391));
NOR2XL cynw_cm_float_cos_I4784 (.Y(N15280), .A(N15541), .B(N14961));
OAI2BB2XL cynw_cm_float_cos_I4785 (.Y(N15424), .A0N(N15455), .A1N(N15276), .B0(N15309), .B1(N15108));
NOR2XL cynw_cm_float_cos_I4786 (.Y(N15575), .A(N15309), .B(N15246));
INVXL cynw_cm_float_cos_I4787 (.Y(N15378), .A(N15096));
INVXL cynw_cm_float_cos_I4788 (.Y(N15530), .A(N15235));
INVXL cynw_cm_float_cos_I4789 (.Y(N15012), .A(N15367));
INVXL cynw_cm_float_cos_I4790 (.Y(N15154), .A(N14999));
AOI21X1 cynw_cm_float_cos_I4791 (.Y(N15550), .A0(N15427), .A1(N15096), .B0(N15281));
AOI21X1 cynw_cm_float_cos_I4792 (.Y(N15175), .A0(N15057), .A1(N15235), .B0(N15578));
AOI21X1 cynw_cm_float_cos_I4793 (.Y(N15463), .A0(N15367), .A1(N15343), .B0(N15200));
AOI21XL cynw_cm_float_cos_I4794 (.Y(N15091), .A0(N14973), .A1(N14999), .B0(N15490));
AOI21X2 cynw_cm_float_cos_I4795 (.Y(N15376), .A0(N15255), .A1(N15281), .B0(N15117));
NAND2X2 cynw_cm_float_cos_I4796 (.Y(N15524), .A(N15255), .B(N15427));
AOI21X1 cynw_cm_float_cos_I4797 (.Y(N15008), .A0(N15554), .A1(N15578), .B0(N15402));
NAND2XL cynw_cm_float_cos_I4798 (.Y(N15152), .A(N15554), .B(N15057));
AOI21X1 cynw_cm_float_cos_I4799 (.Y(N15290), .A0(N15176), .A1(N15200), .B0(N15036));
NAND2XL cynw_cm_float_cos_I4800 (.Y(N15435), .A(N15343), .B(N15176));
AOI21X2 cynw_cm_float_cos_I4801 (.Y(N15587), .A0(N15464), .A1(N15490), .B0(N15320));
NAND2X1 cynw_cm_float_cos_I4802 (.Y(N15064), .A(N15464), .B(N14973));
AOI21X2 cynw_cm_float_cos_I4803 (.Y(N15207), .A0(N15094), .A1(N15117), .B0(N14948));
NAND2X1 cynw_cm_float_cos_I4804 (.Y(N15352), .A(N15094), .B(N15255));
AOI21X2 cynw_cm_float_cos_I4805 (.Y(N15499), .A0(N15377), .A1(N15402), .B0(N15232));
NAND2X1 cynw_cm_float_cos_I4806 (.Y(N14981), .A(N15377), .B(N15554));
AOI21X2 cynw_cm_float_cos_I4807 (.Y(N15127), .A0(N15009), .A1(N15036), .B0(N15528));
NAND2XL cynw_cm_float_cos_I4808 (.Y(N15265), .A(N15009), .B(N15176));
AOI21X2 cynw_cm_float_cos_I4809 (.Y(N15409), .A0(N15295), .A1(N15320), .B0(N15153));
NAND2XL cynw_cm_float_cos_I4810 (.Y(N15565), .A(N15295), .B(N15464));
AOI21X2 cynw_cm_float_cos_I4811 (.Y(N15044), .A0(N15588), .A1(N14948), .B0(N15437));
NAND2X2 cynw_cm_float_cos_I4812 (.Y(N15184), .A(N15588), .B(N15094));
AOI21X1 cynw_cm_float_cos_I4813 (.Y(N15330), .A0(N15208), .A1(N15232), .B0(N15069));
NAND2XL cynw_cm_float_cos_I4814 (.Y(N15473), .A(N15208), .B(N15377));
AOI21X1 cynw_cm_float_cos_I4815 (.Y(N14956), .A0(N15503), .A1(N15528), .B0(N15353));
NAND2XL cynw_cm_float_cos_I4816 (.Y(N15105), .A(N15503), .B(N15009));
AOI21X1 cynw_cm_float_cos_I4817 (.Y(N15241), .A0(N15128), .A1(N15153), .B0(N14982));
NAND2X1 cynw_cm_float_cos_I4818 (.Y(N15386), .A(N15295), .B(N15128));
AOI21XL cynw_cm_float_cos_I4819 (.Y(N15539), .A0(N15410), .A1(N15437), .B0(N15268));
NAND2XL cynw_cm_float_cos_I4820 (.Y(N15019), .A(N15588), .B(N15410));
AOI21X1 cynw_cm_float_cos_I4821 (.Y(N15161), .A0(N15047), .A1(N15069), .B0(N15566));
NAND2X1 cynw_cm_float_cos_I4822 (.Y(N15306), .A(N15208), .B(N15047));
AOI21XL cynw_cm_float_cos_I4823 (.Y(N15448), .A0(N15331), .A1(N15353), .B0(N15185));
NAND2XL cynw_cm_float_cos_I4824 (.Y(N15597), .A(N15331), .B(N15503));
AOI21XL cynw_cm_float_cos_I4825 (.Y(N15081), .A0(N14957), .A1(N14982), .B0(N15477));
NAND2X1 cynw_cm_float_cos_I4826 (.Y(N15219), .A(N14957), .B(N15128));
AOI21XL cynw_cm_float_cos_I4827 (.Y(N15361), .A0(N15244), .A1(N15268), .B0(N15106));
NAND2XL cynw_cm_float_cos_I4828 (.Y(N15513), .A(N15244), .B(N15410));
AOI21XL cynw_cm_float_cos_I4829 (.Y(N14992), .A0(N15540), .A1(N15566), .B0(N15387));
NAND2XL cynw_cm_float_cos_I4830 (.Y(N15135), .A(N15540), .B(N15047));
AOI21XL cynw_cm_float_cos_I4831 (.Y(N15278), .A0(N15162), .A1(N15185), .B0(N15024));
NAND2XL cynw_cm_float_cos_I4832 (.Y(N15420), .A(N15162), .B(N15331));
AOI21XL cynw_cm_float_cos_I4833 (.Y(N15573), .A0(N15451), .A1(N15477), .B0(N15307));
NAND2XL cynw_cm_float_cos_I4834 (.Y(N15054), .A(N15451), .B(N14957));
AOI21XL cynw_cm_float_cos_I4835 (.Y(N15195), .A0(N15082), .A1(N15106), .B0(N15599));
NAND2XL cynw_cm_float_cos_I4836 (.Y(N15338), .A(N15082), .B(N15244));
AOI21XL cynw_cm_float_cos_I4837 (.Y(N15487), .A0(N15363), .A1(N15387), .B0(N15223));
NAND2XL cynw_cm_float_cos_I4838 (.Y(N14967), .A(N15363), .B(N15540));
AOI21XL cynw_cm_float_cos_I4839 (.Y(N15113), .A0(N14997), .A1(N15024), .B0(N15515));
NAND2XL cynw_cm_float_cos_I4840 (.Y(N15253), .A(N14997), .B(N15162));
AOI21XL cynw_cm_float_cos_I4841 (.Y(N15399), .A0(N15280), .A1(N15307), .B0(N15137));
NAND2XL cynw_cm_float_cos_I4842 (.Y(N15547), .A(N15280), .B(N15451));
AOI21XL cynw_cm_float_cos_I4843 (.Y(N15032), .A0(N15575), .A1(N15599), .B0(N15424));
NAND2XL cynw_cm_float_cos_I4844 (.Y(N15172), .A(N15575), .B(N15082));
INVXL cynw_cm_float_cos_I4845 (.Y(N15297), .A(N15378));
INVXL cynw_cm_float_cos_I4846 (.Y(N15441), .A(N15530));
INVXL cynw_cm_float_cos_I4847 (.Y(N15589), .A(N15012));
INVXL cynw_cm_float_cos_I4848 (.Y(N15071), .A(N15154));
INVXL cynw_cm_float_cos_I4849 (.Y(N15211), .A(N15550));
INVXL cynw_cm_float_cos_I4850 (.Y(N15354), .A(N15175));
INVXL cynw_cm_float_cos_I4851 (.Y(N15505), .A(N15463));
INVXL cynw_cm_float_cos_I4852 (.Y(N14985), .A(N15091));
OAI21XL cynw_cm_float_cos_I4853 (.Y(N14978), .A0(N15524), .A1(N15378), .B0(N15376));
OAI21X1 cynw_cm_float_cos_I4854 (.Y(N15261), .A0(N15530), .A1(N15152), .B0(N15008));
OAI21XL cynw_cm_float_cos_I4855 (.Y(N15562), .A0(N15012), .A1(N15435), .B0(N15290));
OAI21X1 cynw_cm_float_cos_I4856 (.Y(N15181), .A0(N15064), .A1(N15154), .B0(N15587));
OAI21X1 cynw_cm_float_cos_I4857 (.Y(N15469), .A0(N15550), .A1(N15352), .B0(N15207));
OAI21XL cynw_cm_float_cos_I4858 (.Y(N15102), .A0(N14981), .A1(N15175), .B0(N15499));
OAI21XL cynw_cm_float_cos_I4859 (.Y(N15383), .A0(N15265), .A1(N15463), .B0(N15127));
OAI21XL cynw_cm_float_cos_I4860 (.Y(N15015), .A0(N15565), .A1(N15091), .B0(N15409));
OAI21X2 cynw_cm_float_cos_I4861 (.Y(N15303), .A0(N15184), .A1(N15376), .B0(N15044));
NOR2X2 cynw_cm_float_cos_I4862 (.Y(N15444), .A(N15184), .B(N15524));
OAI21X1 cynw_cm_float_cos_I4863 (.Y(N15594), .A0(N15473), .A1(N15008), .B0(N15330));
NOR2XL cynw_cm_float_cos_I4864 (.Y(N15078), .A(N15473), .B(N15152));
OAI21XL cynw_cm_float_cos_I4865 (.Y(N15215), .A0(N15105), .A1(N15290), .B0(N14956));
NOR2X1 cynw_cm_float_cos_I4866 (.Y(N15358), .A(N15105), .B(N15435));
OAI21X1 cynw_cm_float_cos_I4867 (.Y(N15510), .A0(N15386), .A1(N15587), .B0(N15241));
NOR2X1 cynw_cm_float_cos_I4868 (.Y(N14988), .A(N15386), .B(N15064));
OAI21X1 cynw_cm_float_cos_I4869 (.Y(N15132), .A0(N15019), .A1(N15207), .B0(N15539));
NOR2XL cynw_cm_float_cos_I4870 (.Y(N15275), .A(N15019), .B(N15352));
OAI21X1 cynw_cm_float_cos_I4871 (.Y(N15416), .A0(N15306), .A1(N15499), .B0(N15161));
NOR2X1 cynw_cm_float_cos_I4872 (.Y(N15571), .A(N15306), .B(N14981));
OAI21XL cynw_cm_float_cos_I4873 (.Y(N15052), .A0(N15597), .A1(N15127), .B0(N15448));
NOR2XL cynw_cm_float_cos_I4874 (.Y(N15190), .A(N15597), .B(N15265));
OAI21X1 cynw_cm_float_cos_I4875 (.Y(N15334), .A0(N15219), .A1(N15409), .B0(N15081));
NOR2X1 cynw_cm_float_cos_I4876 (.Y(N15483), .A(N15219), .B(N15565));
OAI21XL cynw_cm_float_cos_I4877 (.Y(N14963), .A0(N15513), .A1(N15044), .B0(N15361));
NOR2XL cynw_cm_float_cos_I4878 (.Y(N15110), .A(N15513), .B(N15184));
OAI21XL cynw_cm_float_cos_I4879 (.Y(N15249), .A0(N15135), .A1(N15330), .B0(N14992));
NOR2XL cynw_cm_float_cos_I4880 (.Y(N15393), .A(N15135), .B(N15473));
OAI21XL cynw_cm_float_cos_I4881 (.Y(N15543), .A0(N15420), .A1(N14956), .B0(N15278));
NOR2XL cynw_cm_float_cos_I4882 (.Y(N15028), .A(N15420), .B(N15105));
OAI21XL cynw_cm_float_cos_I4883 (.Y(N15166), .A0(N15054), .A1(N15241), .B0(N15573));
NOR2XL cynw_cm_float_cos_I4884 (.Y(N15312), .A(N15054), .B(N15386));
OAI21XL cynw_cm_float_cos_I4885 (.Y(N15457), .A0(N15338), .A1(N15539), .B0(N15195));
NOR2XL cynw_cm_float_cos_I4886 (.Y(N14940), .A(N15338), .B(N15019));
OAI21XL cynw_cm_float_cos_I4887 (.Y(N15086), .A0(N14967), .A1(N15161), .B0(N15487));
NOR2XL cynw_cm_float_cos_I4888 (.Y(N15226), .A(N14967), .B(N15306));
OAI21XL cynw_cm_float_cos_I4889 (.Y(N15369), .A0(N15253), .A1(N15448), .B0(N15113));
NOR2XL cynw_cm_float_cos_I4890 (.Y(N15518), .A(N15253), .B(N15597));
OAI21XL cynw_cm_float_cos_I4891 (.Y(N15001), .A0(N15547), .A1(N15081), .B0(N15399));
NOR2XL cynw_cm_float_cos_I4892 (.Y(N15143), .A(N15547), .B(N15219));
OAI21X1 cynw_cm_float_cos_I4893 (.Y(N15283), .A0(N15172), .A1(N15361), .B0(N15032));
NOR2X1 cynw_cm_float_cos_I4894 (.Y(N15428), .A(N15513), .B(N15172));
INVXL cynw_cm_float_cos_I4895 (.Y(N15412), .A(N15297));
AOI21XL cynw_cm_float_cos_I4896 (.Y(N15567), .A0(N15444), .A1(N15297), .B0(N15303));
AOI21X1 cynw_cm_float_cos_I4897 (.Y(N15187), .A0(N15078), .A1(N15441), .B0(N15594));
AOI21X1 cynw_cm_float_cos_I4898 (.Y(N15479), .A0(N15358), .A1(N15589), .B0(N15215));
AOI21X1 cynw_cm_float_cos_I4899 (.Y(N15107), .A0(N14988), .A1(N15071), .B0(N15510));
AOI21X1 cynw_cm_float_cos_I4900 (.Y(N15390), .A0(N15275), .A1(N15211), .B0(N15132));
AOI21X1 cynw_cm_float_cos_I4901 (.Y(N15026), .A0(N15571), .A1(N15354), .B0(N15416));
AOI21XL cynw_cm_float_cos_I4902 (.Y(N15308), .A0(N15190), .A1(N15505), .B0(N15052));
AOI21X1 cynw_cm_float_cos_I4903 (.Y(N14938), .A0(N15483), .A1(N14985), .B0(N15334));
AOI21X1 cynw_cm_float_cos_I4904 (.Y(N15225), .A0(N15110), .A1(N14978), .B0(N14963));
AOI21XL cynw_cm_float_cos_I4905 (.Y(N15516), .A0(N15393), .A1(N15261), .B0(N15249));
AOI21XL cynw_cm_float_cos_I4906 (.Y(N15140), .A0(N15028), .A1(N15562), .B0(N15543));
AOI21XL cynw_cm_float_cos_I4907 (.Y(N15426), .A0(N15312), .A1(N15181), .B0(N15166));
AOI21X1 cynw_cm_float_cos_I4908 (.Y(N15056), .A0(N14940), .A1(N15469), .B0(N15457));
AOI21XL cynw_cm_float_cos_I4909 (.Y(N15342), .A0(N15226), .A1(N15102), .B0(N15086));
AOI21XL cynw_cm_float_cos_I4910 (.Y(N14972), .A0(N15518), .A1(N15383), .B0(N15369));
AOI21X2 cynw_cm_float_cos_I4911 (.Y(N15553), .A0(N15428), .A1(N15303), .B0(N15283));
NAND2X1 cynw_cm_float_cos_I4912 (.Y(N15035), .A(N15428), .B(N15444));
AO21XL cynw_cm_float_cos_I4913 (.Y(N15366), .A0(N15143), .A1(N15015), .B0(N15001));
OAI21X4 cynw_cm_float_cos_I4914 (.Y(inst_cellmath__201[49]), .A0(N15035), .A1(N15412), .B0(N15553));
NAND2BXL cynw_cm_float_cos_I4923 (.Y(N14991), .AN(N15549), .B(N15034));
NAND2BXL cynw_cm_float_cos_I4924 (.Y(N15419), .AN(N15173), .B(N15317));
NAND2BXL cynw_cm_float_cos_I4925 (.Y(N15192), .AN(N15462), .B(N14946));
NAND2BXL cynw_cm_float_cos_I4926 (.Y(N14966), .AN(N15090), .B(N15231));
NAND2BXL cynw_cm_float_cos_I4927 (.Y(N15397), .AN(N15374), .B(N15523));
NAND2BXL cynw_cm_float_cos_I4928 (.Y(N15170), .AN(N15007), .B(N15150));
NAND2BXL cynw_cm_float_cos_I4929 (.Y(N14944), .AN(N15289), .B(N15434));
NAND2BXL cynw_cm_float_cos_I4930 (.Y(N15372), .AN(N15585), .B(N15063));
NAND2BXL cynw_cm_float_cos_I4931 (.Y(N15147), .AN(N15206), .B(N15350));
NAND2BXL cynw_cm_float_cos_I4932 (.Y(N15583), .AN(N15496), .B(N14980));
NAND2BXL cynw_cm_float_cos_I4933 (.Y(N15348), .AN(N15125), .B(N15263));
NAND2BXL cynw_cm_float_cos_I4934 (.Y(N15123), .AN(N15408), .B(N15563));
NAND2BXL cynw_cm_float_cos_I4935 (.Y(N15559), .AN(N15042), .B(N15183));
NAND2BXL cynw_cm_float_cos_I4936 (.Y(N15325), .AN(N15328), .B(N15471));
NAND2BXL cynw_cm_float_cos_I4937 (.Y(N15100), .AN(N14955), .B(N15103));
NAND2BXL cynw_cm_float_cos_I4938 (.Y(N15534), .AN(N15239), .B(N15385));
NAND2BXL cynw_cm_float_cos_I4939 (.Y(N15301), .AN(N15536), .B(N15017));
NAND2BXL cynw_cm_float_cos_I4940 (.Y(N15075), .AN(N15160), .B(N15304));
NAND2BXL cynw_cm_float_cos_I4941 (.Y(N15508), .AN(N15446), .B(N15596));
NAND2BXL cynw_cm_float_cos_I4942 (.Y(N15273), .AN(N15079), .B(N15217));
NAND2BXL cynw_cm_float_cos_I4943 (.Y(N15050), .AN(N15360), .B(N15511));
NAND2BXL cynw_cm_float_cos_I4944 (.Y(N15481), .AN(N14990), .B(N15134));
NAND2BXL cynw_cm_float_cos_I4945 (.Y(N15247), .AN(N15276), .B(N15418));
XOR2XL cynw_cm_float_cos_I4954 (.Y(inst_cellmath__201[25]), .A(N14978), .B(N14991));
XOR2XL cynw_cm_float_cos_I4955 (.Y(inst_cellmath__201[26]), .A(N15261), .B(N15419));
XOR2XL cynw_cm_float_cos_I4956 (.Y(inst_cellmath__201[27]), .A(N15562), .B(N15192));
XOR2XL cynw_cm_float_cos_I4957 (.Y(inst_cellmath__201[28]), .A(N15181), .B(N14966));
XOR2XL cynw_cm_float_cos_I4958 (.Y(inst_cellmath__201[29]), .A(N15469), .B(N15397));
XOR2XL cynw_cm_float_cos_I4959 (.Y(inst_cellmath__201[30]), .A(N15102), .B(N15170));
XOR2XL cynw_cm_float_cos_I4960 (.Y(inst_cellmath__201[31]), .A(N15383), .B(N14944));
XOR2XL cynw_cm_float_cos_I4961 (.Y(inst_cellmath__201[32]), .A(N15372), .B(N15015));
INVXL xnor2_A_I11478 (.Y(N23433), .A(N15567));
MXI2XL xnor2_A_I11479 (.Y(inst_cellmath__201[33]), .A(N15567), .B(N23433), .S0(N15147));
XNOR2XL cynw_cm_float_cos_I4963 (.Y(inst_cellmath__201[34]), .A(N15583), .B(N15187));
INVXL xnor2_A_I11480 (.Y(N23439), .A(N15479));
MXI2XL xnor2_A_I11481 (.Y(inst_cellmath__201[35]), .A(N15479), .B(N23439), .S0(N15348));
XNOR2XL cynw_cm_float_cos_I4965 (.Y(inst_cellmath__201[36]), .A(N15123), .B(N15107));
XNOR2XL cynw_cm_float_cos_I4966 (.Y(inst_cellmath__201[37]), .A(N15559), .B(N15390));
XNOR2XL cynw_cm_float_cos_I4967 (.Y(inst_cellmath__201[38]), .A(N15325), .B(N15026));
XNOR2XL cynw_cm_float_cos_I4968 (.Y(inst_cellmath__201[39]), .A(N15100), .B(N15308));
INVXL xnor2_A_I30589 (.Y(N45805), .A(N14938));
MXI2XL xnor2_A_I30590 (.Y(inst_cellmath__201[40]), .A(N14938), .B(N45805), .S0(N15534));
INVXL xnor2_A_I30591 (.Y(N45811), .A(N15301));
MXI2XL xnor2_A_I30592 (.Y(inst_cellmath__201[41]), .A(N15301), .B(N45811), .S0(N15225));
INVXL xnor2_A_I30593 (.Y(N45817), .A(N15075));
MXI2XL xnor2_A_I30594 (.Y(inst_cellmath__201[42]), .A(N15075), .B(N45817), .S0(N15516));
INVXL xnor2_A_I30595 (.Y(N45823), .A(N15508));
MXI2XL xnor2_A_I30596 (.Y(inst_cellmath__201[43]), .A(N15508), .B(N45823), .S0(N15140));
INVXL xnor2_A_I30597 (.Y(N45829), .A(N15273));
MXI2XL xnor2_A_I30598 (.Y(inst_cellmath__201[44]), .A(N15273), .B(N45829), .S0(N15426));
INVXL xnor2_A_I30599 (.Y(N45835), .A(N15050));
MXI2XL xnor2_A_I30600 (.Y(inst_cellmath__201[45]), .A(N15050), .B(N45835), .S0(N15056));
INVXL xnor2_A_I30601 (.Y(N45841), .A(N15481));
MXI2XL xnor2_A_I30602 (.Y(inst_cellmath__201[46]), .A(N15481), .B(N45841), .S0(N15342));
INVXL xnor2_A_I30603 (.Y(N45847), .A(N15247));
MXI2XL xnor2_A_I30604 (.Y(inst_cellmath__201[47]), .A(N15247), .B(N45847), .S0(N14972));
INVX6 inst_cellmath__200_0_I4978 (.Y(N16220), .A(inst_cellmath__201[49]));
AND2XL inst_cellmath__200_0_I5004 (.Y(inst_cellmath__210[0]), .A(inst_cellmath__201[25]), .B(N16220));
AND2X1 inst_cellmath__200_0_I5005 (.Y(inst_cellmath__210[1]), .A(N16220), .B(inst_cellmath__201[26]));
AND2XL inst_cellmath__200_0_I5006 (.Y(inst_cellmath__210[2]), .A(inst_cellmath__201[27]), .B(N16220));
CLKAND2X2 inst_cellmath__200_0_I5007 (.Y(inst_cellmath__210[3]), .A(inst_cellmath__201[28]), .B(N16220));
CLKAND2X3 inst_cellmath__200_0_I5008 (.Y(inst_cellmath__210[4]), .A(inst_cellmath__201[29]), .B(N16220));
AND2X1 inst_cellmath__200_0_I5009 (.Y(inst_cellmath__210[5]), .A(N16220), .B(inst_cellmath__201[30]));
AND2X1 inst_cellmath__200_0_I5010 (.Y(inst_cellmath__210[6]), .A(N16220), .B(inst_cellmath__201[31]));
CLKAND2X2 inst_cellmath__200_0_I5011 (.Y(inst_cellmath__210[7]), .A(inst_cellmath__201[32]), .B(N16220));
CLKAND2X2 inst_cellmath__200_0_I5012 (.Y(inst_cellmath__210[8]), .A(N16220), .B(inst_cellmath__201[33]));
CLKAND2X2 inst_cellmath__200_0_I5013 (.Y(inst_cellmath__210[9]), .A(inst_cellmath__201[34]), .B(N16220));
CLKAND2X2 inst_cellmath__200_0_I5014 (.Y(inst_cellmath__210[10]), .A(N16220), .B(inst_cellmath__201[35]));
NAND2X1 inst_cellmath__200_0_I10417 (.Y(N23255), .A(inst_cellmath__201[36]), .B(N16220));
INVX2 inst_cellmath__200_0_I10418 (.Y(inst_cellmath__210[11]), .A(N23255));
NAND2X1 inst_cellmath__200_0_I10643 (.Y(N23324), .A(inst_cellmath__201[37]), .B(N16220));
INVX1 inst_cellmath__200_0_I10644 (.Y(inst_cellmath__210[12]), .A(N23324));
CLKAND2X2 inst_cellmath__200_0_I5017 (.Y(inst_cellmath__210[13]), .A(inst_cellmath__201[38]), .B(N16220));
NAND2X1 inst_cellmath__200_0_I10655 (.Y(N23358), .A(inst_cellmath__201[39]), .B(N16220));
INVX2 inst_cellmath__200_0_I10656 (.Y(inst_cellmath__210[14]), .A(N23358));
AND2XL inst_cellmath__200_0_I5019 (.Y(inst_cellmath__210[15]), .A(inst_cellmath__201[40]), .B(N16220));
AND2X1 inst_cellmath__200_0_I5020 (.Y(inst_cellmath__210[16]), .A(N16220), .B(inst_cellmath__201[41]));
AND2X1 inst_cellmath__200_0_I5021 (.Y(inst_cellmath__210[17]), .A(N16220), .B(inst_cellmath__201[42]));
AND2X1 inst_cellmath__200_0_I5022 (.Y(inst_cellmath__210[18]), .A(N16220), .B(inst_cellmath__201[43]));
AND2X1 inst_cellmath__200_0_I5023 (.Y(inst_cellmath__210[19]), .A(N16220), .B(inst_cellmath__201[44]));
AND2X1 inst_cellmath__200_0_I10629 (.Y(inst_cellmath__210[20]), .A(N16220), .B(inst_cellmath__201[45]));
AND2X1 inst_cellmath__200_0_I5025 (.Y(inst_cellmath__210[21]), .A(N16220), .B(inst_cellmath__201[46]));
AND2X1 inst_cellmath__200_0_I5026 (.Y(inst_cellmath__210[22]), .A(inst_cellmath__201[47]), .B(N16220));
OR4X1 inst_cellmath__17_0_I30037 (.Y(N16294), .A(a_exp[7]), .B(a_exp[6]), .C(a_exp[0]), .D(a_exp[5]));
OR4X1 inst_cellmath__17_0_I30038 (.Y(N16298), .A(a_exp[4]), .B(a_exp[2]), .C(a_exp[3]), .D(a_exp[1]));
NAND2XL inst_cellmath__21_0_I5038 (.Y(N16328), .A(a_exp[2]), .B(a_exp[1]));
NOR2XL inst_cellmath__21_0_I5039 (.Y(N16334), .A(a_exp[3]), .B(a_exp[4]));
NAND2XL inst_cellmath__21_0_I5040 (.Y(N16332), .A(a_exp[5]), .B(a_exp[6]));
AOI21XL inst_cellmath__21_0_I5041 (.Y(N16324), .A0(N16328), .A1(N16334), .B0(N16332));
NAND2XL inst_cellmath__19_0_I5048 (.Y(N16362), .A(a_exp[4]), .B(a_exp[3]));
NOR2XL inst_cellmath__19_0_I5051 (.Y(N16357), .A(N16362), .B(N16328));
NOR2XL inst_cellmath__19_0_I29502 (.Y(inst_cellmath__42[8]), .A(N7291), .B(N7267));
XOR2XL inst_cellmath__19_0_I29503 (.Y(N45155), .A(N15366), .B(N15455));
NAND2XL inst_cellmath__19_0_I29504 (.Y(N45117), .A(inst_cellmath__61[22]), .B(N16220));
NOR2XL inst_cellmath__19_0_I29505 (.Y(N45128), .A(inst_cellmath__42[7]), .B(inst_cellmath__42[6]));
OA22X1 inst_cellmath__19_0_I30039 (.Y(N45139), .A0(a_exp[7]), .A1(N16324), .B0(N16294), .B1(N16298));
NAND2XL inst_cellmath__19_0_I29507 (.Y(N45150), .A(a_exp[6]), .B(a_exp[5]));
NAND3XL inst_cellmath__19_0_I29509 (.Y(N45152), .A(a_exp[7]), .B(a_exp[0]), .C(N16357));
NOR2XL inst_cellmath__19_0_I29510 (.Y(inst_cellmath__19), .A(N45150), .B(N45152));
NAND2XL cynw_cm_float_cos_I5083 (.Y(N16464), .A(a_sign), .B(inst_cellmath__19));
NOR2XL inst_cellmath__24_0_I5060 (.Y(N16380), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__24_0_I5061 (.Y(N16390), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__24_0_I5062 (.Y(N16401), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__24_0_I5063 (.Y(N16411), .A(a_man[4]), .B(a_man[3]));
AND4XL inst_cellmath__24_0_I30042 (.Y(N16393), .A(N16411), .B(N16380), .C(N16390), .D(N16401));
NOR2XL inst_cellmath__24_0_I5055 (.Y(N16376), .A(a_man[20]), .B(a_man[19]));
NOR2XL inst_cellmath__24_0_I5053 (.Y(N16403), .A(a_man[0]), .B(a_man[1]));
NOR2XL inst_cellmath__24_0_I5056 (.Y(N16386), .A(a_man[18]), .B(a_man[17]));
NOR2XL inst_cellmath__24_0_I5057 (.Y(N16397), .A(a_man[16]), .B(a_man[15]));
NOR2XL inst_cellmath__24_0_I5058 (.Y(N16407), .A(a_man[14]), .B(a_man[13]));
NOR2XL inst_cellmath__24_0_I5059 (.Y(N16417), .A(a_man[12]), .B(a_man[11]));
AND4XL inst_cellmath__24_0_I30045 (.Y(N16409), .A(N16417), .B(N16386), .C(N16397), .D(N16407));
NAND3XL inst_cellmath__24_0_I11484 (.Y(N23456), .A(N6122), .B(N16403), .C(N16409));
NAND4BXL inst_cellmath__24_0_I30047 (.Y(inst_cellmath__24), .AN(N23456), .B(N6213), .C(N16393), .D(N16376));
NOR2XL inst_cellmath__19_0_I29508 (.Y(N45159), .A(N16464), .B(inst_cellmath__24));
NOR3BXL inst_cellmath__19_0_I29511 (.Y(N45122), .AN(inst_cellmath__19), .B(a_sign), .C(inst_cellmath__24));
NOR2XL inst_cellmath__19_0_I29512 (.Y(N45119), .A(N45122), .B(N45159));
OR2XL inst_cellmath__19_0_I29513 (.Y(inst_cellmath__68), .A(N45159), .B(N45122));
NOR2X2 inst_cellmath__211__182__I5120 (.Y(N16550), .A(inst_cellmath__210[22]), .B(inst_cellmath__210[21]));
NOR2X1 inst_cellmath__211__182__I5119 (.Y(N16531), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[19]));
NAND2X1 inst_cellmath__211__182__I5134 (.Y(N16528), .A(N16531), .B(N16550));
NOR2X1 inst_cellmath__211__182__I5116 (.Y(N16523), .A(inst_cellmath__210[17]), .B(inst_cellmath__210[18]));
NOR2X1 inst_cellmath__211__182__I5115 (.Y(N16505), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[15]));
NAND2X1 inst_cellmath__211__182__I5133 (.Y(N16511), .A(N16505), .B(N16523));
NOR2X2 inst_cellmath__211__182__I5140 (.Y(N16544), .A(N16528), .B(N16511));
NOR2X4 inst_cellmath__211__182__I5105 (.Y(N16558), .A(inst_cellmath__210[9]), .B(inst_cellmath__210[10]));
NOR2X4 inst_cellmath__211__182__I5104 (.Y(N16538), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]));
NAND2X4 inst_cellmath__211__182__I5128 (.Y(N16571), .A(N16538), .B(N16558));
NOR2X2 inst_cellmath__211__182__I5099 (.Y(N16529), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[5]));
NOR2X2 inst_cellmath__211__182__I5098 (.Y(N16512), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[3]));
NAND2X2 inst_cellmath__211__182__I5124 (.Y(N16565), .A(N16529), .B(N16512));
INVXL inst_cellmath__211__182__I5135 (.Y(N16508), .A(N16565));
NOR2X4 inst_cellmath__211__182__I5111 (.Y(N16498), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[13]));
NOR2X2 inst_cellmath__211__182__I5110 (.Y(N16567), .A(inst_cellmath__210[11]), .B(inst_cellmath__210[12]));
NAND2X4 inst_cellmath__211__182__I5129 (.Y(N16503), .A(N16498), .B(N16567));
INVXL inst_cellmath__211__182__I5136 (.Y(N16545), .A(N16503));
OAI21XL inst_cellmath__211__182__I5137 (.Y(N16566), .A0(N16571), .A1(N16508), .B0(N16545));
NAND2BXL inst_cellmath__211__182__I5139 (.Y(N16504), .AN(N16528), .B(N16511));
INVX2 inst_cellmath__220__188__I29674 (.Y(N16494), .A(N16544));
OAI21X1 inst_cellmath__211__182__I5144 (.Y(N550), .A0(N16566), .A1(N16494), .B0(N16504));
NOR2X4 inst_cellmath__211__182__I5138 (.Y(N16517), .A(N16503), .B(N16571));
OR2XL inst_cellmath__211__182__I5121 (.Y(N16556), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[1]));
INVXL inst_cellmath__211__182__I5122 (.Y(N16506), .A(N16529));
AOI21XL inst_cellmath__211__182__I5123 (.Y(N16525), .A0(N16512), .A1(N16556), .B0(N16506));
NAND2BXL inst_cellmath__211__182__I5125 (.Y(N16515), .AN(N16538), .B(N16558));
INVXL inst_cellmath__211__182__I5126 (.Y(N16533), .A(N16498));
AOI21X1 inst_cellmath__211__182__I5127 (.Y(N16551), .A0(N16567), .A1(N16515), .B0(N16533));
NAND2BXL inst_cellmath__211__182__I5130 (.Y(N16541), .AN(N16505), .B(N16523));
INVXL inst_cellmath__211__182__I5131 (.Y(N16561), .A(N16550));
AOI21XL inst_cellmath__211__182__I5132 (.Y(N16492), .A0(N16531), .A1(N16541), .B0(N16561));
INVXL inst_cellmath__211__182__I5091 (.Y(N16497), .A(inst_cellmath__210[0]));
INVXL inst_cellmath__211__182__I5092 (.Y(N16534), .A(inst_cellmath__210[2]));
OAI21X2 inst_cellmath__211__182__I5093 (.Y(N16552), .A0(inst_cellmath__210[1]), .A1(N16497), .B0(N16534));
INVX3 inst_cellmath__211__182__I5094 (.Y(N16522), .A(inst_cellmath__210[3]));
NOR2X4 inst_cellmath__211__182__I5095 (.Y(N16542), .A(inst_cellmath__210[4]), .B(N16522));
INVX1 inst_cellmath__211__182__I5096 (.Y(N16562), .A(inst_cellmath__210[6]));
OAI21X2 inst_cellmath__211__182__I5097 (.Y(N16493), .A0(inst_cellmath__210[5]), .A1(N16542), .B0(N16562));
OAI21X2 inst_cellmath__211__182__I5148 (.Y(N16537), .A0(N16565), .A1(N16552), .B0(N16493));
INVX2 inst_cellmath__211__182__I5100 (.Y(N16548), .A(inst_cellmath__210[7]));
NOR2X2 inst_cellmath__211__182__I5101 (.Y(N16569), .A(inst_cellmath__210[8]), .B(N16548));
INVXL inst_cellmath__211__182__I5102 (.Y(N16500), .A(inst_cellmath__210[10]));
OAI21X2 inst_cellmath__211__182__I5103 (.Y(N16519), .A0(inst_cellmath__210[9]), .A1(N16569), .B0(N16500));
INVX1 inst_cellmath__211__182__I5106 (.Y(N16489), .A(inst_cellmath__210[11]));
NOR2X2 inst_cellmath__211__182__I5107 (.Y(N16509), .A(inst_cellmath__210[12]), .B(N16489));
INVX1 inst_cellmath__211__182__I5108 (.Y(N16526), .A(inst_cellmath__210[14]));
OAI21X2 inst_cellmath__211__182__I5109 (.Y(N16546), .A0(inst_cellmath__210[13]), .A1(N16509), .B0(N16526));
OAI21X2 inst_cellmath__211__182__I5149 (.Y(N16488), .A0(N16503), .A1(N16519), .B0(N16546));
AOI21X2 inst_cellmath__211__182__I5150 (.Y(N16516), .A0(N16517), .A1(N16537), .B0(N16488));
NOR2BXL inst_cellmath__211__182__I5112 (.Y(N16535), .AN(inst_cellmath__210[15]), .B(inst_cellmath__210[16]));
INVXL inst_cellmath__211__182__I5113 (.Y(N16554), .A(inst_cellmath__210[18]));
OAI21XL inst_cellmath__211__182__I5114 (.Y(N16486), .A0(inst_cellmath__210[17]), .A1(N16535), .B0(N16554));
NOR2BX1 inst_cellmath__211__182__I5117 (.Y(N16564), .AN(inst_cellmath__210[19]), .B(inst_cellmath__210[20]));
INVXL inst_cellmath__211__182__I5090 (.Y(N16557), .A(inst_cellmath__210[22]));
OAI21X1 inst_cellmath__211__182__I5118 (.Y(N16514), .A0(inst_cellmath__210[21]), .A1(N16564), .B0(N16557));
OA21X1 inst_cellmath__211__182__I5151 (.Y(N16553), .A0(N16528), .A1(N16486), .B0(N16514));
AOI21X1 inst_cellmath__220__188__I29675 (.Y(N45547), .A0(N16525), .A1(N16517), .B0(N16551));
INVXL inst_cellmath__220__188__I29676 (.Y(N45552), .A(N16492));
OAI21X1 inst_cellmath__220__188__I29677 (.Y(N549), .A0(N16494), .A1(N45547), .B0(N45552));
OAI21X2 inst_cellmath__220__188__I29678 (.Y(N548), .A0(N16494), .A1(N16516), .B0(N16553));
AND2XL cynw_cm_float_cos_I5154 (.Y(N16636), .A(N548), .B(N549));
NAND2BXL inst_cellmath__220__188__I29453 (.Y(N551), .AN(N16517), .B(N16544));
INVXL gen2_alt_A_I30605 (.Y(N45854), .A(N551));
OAI2BB1X1 gen2_alt_A_I30606 (.Y(N16646), .A0N(N16636), .A1N(N550), .B0(N45854));
XNOR2X1 cynw_cm_float_cos_I10811 (.Y(inst_cellmath__215[4]), .A(N16494), .B(N16646));
INVX1 inst_cellmath__220__188__I5244 (.Y(N16754), .A(inst_cellmath__215[4]));
INVX3 inst_cellmath__220__188__I5245 (.Y(N16800), .A(N16754));
INVX2 inst_cellmath__220__188__I29679 (.Y(inst_cellmath__215[0]), .A(N548));
INVX3 inst_cellmath__220__188__I5165 (.Y(N16722), .A(inst_cellmath__215[0]));
MX2XL inst_cellmath__220__188__I5176 (.Y(N16694), .A(inst_cellmath__210[8]), .B(inst_cellmath__210[9]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5178 (.Y(N16764), .A(inst_cellmath__210[10]), .B(inst_cellmath__210[11]), .S0(N16722));
XNOR2X1 inst_cellmath__220__188__I29680 (.Y(N45549), .A(N549), .B(inst_cellmath__215[0]));
CLKINVX6 inst_cellmath__220__188__I29681 (.Y(N16759), .A(N45549));
MXI2XL inst_cellmath__220__188__I5202 (.Y(N16815), .A(N16694), .B(N16764), .S0(N16759));
MX2XL inst_cellmath__220__188__I5168 (.Y(N16734), .A(inst_cellmath__210[0]), .B(inst_cellmath__210[1]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5170 (.Y(N16802), .A(inst_cellmath__210[2]), .B(inst_cellmath__210[3]), .S0(N16722));
MXI2XL inst_cellmath__220__188__I5194 (.Y(N16698), .A(N16734), .B(N16802), .S0(N16759));
INVXL inst_cellmath__220__188__I29455 (.Y(N45000), .A(N551));
NAND2XL cynw_cm_float_cos_I5155 (.Y(N16643), .A(N549), .B(N550));
NOR2XL inst_cellmath__220__188__I29454 (.Y(N45002), .A(N16643), .B(inst_cellmath__215[0]));
XNOR2X1 inst_cellmath__220__188__I29458 (.Y(N23318), .A(N45000), .B(N45002));
INVX1 inst_cellmath__220__188__I10614 (.Y(N23319), .A(N23318));
MXI2XL inst_cellmath__220__188__I5231 (.Y(N16762), .A(N16815), .B(N16698), .S0(N23319));
NAND2XL inst_cellmath__19_0_I29514 (.Y(N16808), .A(N16800), .B(N16762));
MX2XL inst_cellmath__220__188__I5180 (.Y(N16669), .A(inst_cellmath__210[12]), .B(inst_cellmath__210[13]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5182 (.Y(N16743), .A(inst_cellmath__210[14]), .B(inst_cellmath__210[15]), .S0(N16722));
MXI2XL inst_cellmath__220__188__I5206 (.Y(N16795), .A(N16669), .B(N16743), .S0(N16759));
MX2XL inst_cellmath__220__188__I5172 (.Y(N16710), .A(inst_cellmath__210[4]), .B(inst_cellmath__210[5]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5174 (.Y(N16782), .A(inst_cellmath__210[6]), .B(inst_cellmath__210[7]), .S0(N16722));
MXI2XL inst_cellmath__220__188__I5198 (.Y(N16675), .A(N16710), .B(N16782), .S0(N16759));
INVX1 inst_cellmath__220__188__I10616 (.Y(N23321), .A(N23318));
MXI2XL inst_cellmath__220__188__I5235 (.Y(N16741), .A(N16795), .B(N16675), .S0(N23321));
NAND2XL inst_cellmath__19_0_I29515 (.Y(N16770), .A(N16741), .B(N16800));
XNOR2X1 cynw_cm_float_cos_I5160 (.Y(inst_cellmath__215[2]), .A(N16636), .B(N550));
CLKINVX6 inst_cellmath__19_0_I29516 (.Y(N16725), .A(inst_cellmath__215[2]));
MXI2XL inst_cellmath__19_0_I30055 (.Y(N45115), .A(N16770), .B(N16808), .S0(N16725));
INVXL inst_cellmath__19_0_I29519 (.Y(N17163), .A(inst_cellmath__19));
NOR2X1 inst_cellmath__19_0_I29520 (.Y(N16991), .A(N45117), .B(N45155));
NAND2BXL inst_cellmath__19_0_I29521 (.Y(N45148), .AN(N16991), .B(N45115));
NOR2XL inst_cellmath__19_0_I29522 (.Y(N45146), .A(inst_cellmath__42[8]), .B(N45128));
OAI21XL inst_cellmath__19_0_I29523 (.Y(N16343), .A0(inst_cellmath__42[8]), .A1(N45128), .B0(N45139));
INVXL inst_cellmath__19_0_I29524 (.Y(N45132), .A(N45139));
NAND2XL inst_cellmath__19_0_I29525 (.Y(N45118), .A(N17163), .B(N45119));
OR3XL inst_cellmath__19_0_I29526 (.Y(N741), .A(N45146), .B(N45132), .C(N45118));
MXI2XL inst_cellmath__19_0_I29527 (.Y(x[15]), .A(N45148), .B(N17163), .S0(N741));
AND2XL inst_cellmath__220__188__I5167 (.Y(N16823), .A(N16722), .B(inst_cellmath__210[0]));
MX2XL inst_cellmath__220__188__I5169 (.Y(N16769), .A(inst_cellmath__210[1]), .B(inst_cellmath__210[2]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5171 (.Y(N16677), .A(inst_cellmath__210[3]), .B(inst_cellmath__210[4]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5173 (.Y(N16749), .A(inst_cellmath__210[5]), .B(inst_cellmath__210[6]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5175 (.Y(N16816), .A(inst_cellmath__210[7]), .B(inst_cellmath__210[8]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5177 (.Y(N16728), .A(inst_cellmath__210[9]), .B(inst_cellmath__210[10]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5179 (.Y(N16796), .A(inst_cellmath__210[11]), .B(inst_cellmath__210[12]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5181 (.Y(N16705), .A(inst_cellmath__210[13]), .B(inst_cellmath__210[14]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5183 (.Y(N16777), .A(inst_cellmath__210[15]), .B(inst_cellmath__210[16]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5184 (.Y(N16811), .A(inst_cellmath__210[16]), .B(inst_cellmath__210[17]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5185 (.Y(N16686), .A(inst_cellmath__210[17]), .B(inst_cellmath__210[18]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5186 (.Y(N16720), .A(inst_cellmath__210[18]), .B(inst_cellmath__210[19]), .S0(N16722));
INVXL inst_cellmath__220__188__I10412 (.Y(N23240), .A(inst_cellmath__210[20]));
NAND2XL inst_cellmath__220__188__I10414 (.Y(N23239), .A(N23240), .B(N16722));
OA21XL inst_cellmath__220__188__I11289 (.Y(N16757), .A0(N16722), .A1(inst_cellmath__210[19]), .B0(N23239));
MX2XL inst_cellmath__220__188__I5188 (.Y(N16790), .A(inst_cellmath__210[20]), .B(inst_cellmath__210[21]), .S0(N16722));
MX2XL inst_cellmath__220__188__I5189 (.Y(N16663), .A(inst_cellmath__210[21]), .B(inst_cellmath__210[22]), .S0(N16722));
NAND2XL inst_cellmath__220__188__I5191 (.Y(N16682), .A(N16823), .B(N16759));
NAND2XL inst_cellmath__220__188__I5192 (.Y(N16755), .A(N16734), .B(N16759));
MXI2X1 inst_cellmath__220__188__I5193 (.Y(N16822), .A(N16823), .B(N16769), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5195 (.Y(N16733), .A(N16769), .B(N16677), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5196 (.Y(N16768), .A(N16802), .B(N16710), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5197 (.Y(N16801), .A(N16677), .B(N16749), .S0(N16759));
MXI2X1 inst_cellmath__220__188__I5199 (.Y(N16709), .A(N16749), .B(N16816), .S0(N16759));
MXI2X1 inst_cellmath__220__188__I5200 (.Y(N16748), .A(N16782), .B(N16694), .S0(N16759));
MXI2X1 inst_cellmath__220__188__I5201 (.Y(N16781), .A(N16816), .B(N16728), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5203 (.Y(N16692), .A(N16728), .B(N16796), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5204 (.Y(N16726), .A(N16764), .B(N16669), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5205 (.Y(N16763), .A(N16796), .B(N16705), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5207 (.Y(N16668), .A(N16705), .B(N16777), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5208 (.Y(N16704), .A(N16743), .B(N16811), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5209 (.Y(N16742), .A(N16777), .B(N16686), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5210 (.Y(N16776), .A(N16811), .B(N16720), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5211 (.Y(N16810), .A(N16686), .B(N16757), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5212 (.Y(N16685), .A(N16720), .B(N16790), .S0(N16759));
MXI2XL inst_cellmath__220__188__I5213 (.Y(N16719), .A(N16757), .B(N16663), .S0(N16759));
XOR2XL inst_cellmath__220__188__I29456 (.Y(inst_cellmath__215[3]), .A(N45002), .B(N551));
INVXL inst_cellmath__220__188__I29457 (.Y(N16681), .A(inst_cellmath__215[3]));
INVX1 inst_cellmath__220__188__I10617 (.Y(N23322), .A(N23318));
INVX2 inst_cellmath__220__188__I10615 (.Y(N23320), .A(N23318));
NOR2XL inst_cellmath__220__188__I5220 (.Y(N16737), .A(N16682), .B(N16681));
NOR2BX1 inst_cellmath__220__188__I30059 (.Y(N16805), .AN(N23318), .B(N16755));
NOR2XL inst_cellmath__220__188__I5222 (.Y(N16715), .A(N16822), .B(N23322));
NOR2XL inst_cellmath__220__188__I5223 (.Y(N16786), .A(N16698), .B(N23321));
NOR2XL inst_cellmath__220__188__I5224 (.Y(N16697), .A(N16733), .B(N23321));
NOR2XL inst_cellmath__220__188__I5225 (.Y(N16767), .A(N16768), .B(N23321));
NOR2XL inst_cellmath__220__188__I5226 (.Y(N16673), .A(N16801), .B(N23321));
NOR2XL inst_cellmath__220__188__I5227 (.Y(N16746), .A(N16675), .B(N23319));
MXI2XL inst_cellmath__220__188__I5228 (.Y(N16814), .A(N16709), .B(N16682), .S0(N23319));
MXI2XL inst_cellmath__220__188__I5229 (.Y(N16691), .A(N16748), .B(N16755), .S0(N23319));
MXI2XL inst_cellmath__220__188__I5230 (.Y(N16724), .A(N16781), .B(N16822), .S0(N23319));
MXI2XL inst_cellmath__220__188__I5232 (.Y(N16794), .A(N16692), .B(N16733), .S0(N16681));
MXI2XL inst_cellmath__220__188__I5233 (.Y(N16667), .A(N16726), .B(N16768), .S0(N23320));
MXI2XL inst_cellmath__220__188__I5234 (.Y(N16703), .A(N16763), .B(N16801), .S0(N23320));
MXI2X1 inst_cellmath__220__188__I5236 (.Y(N16775), .A(N16668), .B(N16709), .S0(N23320));
MXI2X1 inst_cellmath__220__188__I5237 (.Y(N16809), .A(N16704), .B(N16748), .S0(N23320));
MXI2X1 inst_cellmath__220__188__I5238 (.Y(N16684), .A(N16742), .B(N16781), .S0(N23320));
MXI2XL inst_cellmath__220__188__I5239 (.Y(N16718), .A(N16776), .B(N16815), .S0(N23322));
MXI2XL inst_cellmath__220__188__I5240 (.Y(N16756), .A(N16810), .B(N16692), .S0(N23322));
MXI2XL inst_cellmath__220__188__I5241 (.Y(N16789), .A(N16685), .B(N16726), .S0(N23322));
MXI2XL inst_cellmath__220__188__I5242 (.Y(N16662), .A(N16719), .B(N16763), .S0(N23322));
NAND2XL inst_cellmath__220__188__I5249 (.Y(N16680), .A(N16737), .B(N16800));
NAND2XL inst_cellmath__220__188__I5250 (.Y(N16752), .A(N16805), .B(N16800));
NAND2XL inst_cellmath__220__188__I5251 (.Y(N16820), .A(N16715), .B(N16800));
NAND2XL inst_cellmath__220__188__I5252 (.Y(N16731), .A(N16800), .B(N16786));
NAND2XL inst_cellmath__220__188__I5253 (.Y(N16798), .A(N16800), .B(N16697));
NAND2XL inst_cellmath__220__188__I5254 (.Y(N16708), .A(N16800), .B(N16767));
NAND2XL inst_cellmath__220__188__I5255 (.Y(N16780), .A(N16800), .B(N16673));
NAND2XL inst_cellmath__220__188__I5256 (.Y(N16689), .A(N16746), .B(N16800));
NAND2XL inst_cellmath__220__188__I5257 (.Y(N16761), .A(N16814), .B(N16800));
NAND2X1 inst_cellmath__220__188__I5258 (.Y(N16666), .A(N16691), .B(N16800));
NAND2XL inst_cellmath__220__188__I5259 (.Y(N16739), .A(N16724), .B(N16800));
NAND2XL inst_cellmath__220__188__I5261 (.Y(N16717), .A(N16794), .B(N16800));
NAND2X1 inst_cellmath__220__188__I5262 (.Y(N16788), .A(N16667), .B(N16800));
NAND2XL inst_cellmath__220__188__I5263 (.Y(N16699), .A(N16703), .B(N16800));
MXI2X1 inst_cellmath__220__188__I5265 (.Y(N16676), .A(N16737), .B(N16775), .S0(N16800));
MXI2X1 inst_cellmath__220__188__I5266 (.Y(N16711), .A(N16805), .B(N16809), .S0(N16800));
MXI2X1 inst_cellmath__220__188__I5267 (.Y(N16750), .A(N16715), .B(N16684), .S0(N16800));
MXI2XL inst_cellmath__220__188__I5268 (.Y(N16783), .A(N16786), .B(N16718), .S0(N16800));
MXI2XL inst_cellmath__220__188__I5269 (.Y(N16817), .A(N16697), .B(N16756), .S0(N16800));
MXI2XL inst_cellmath__220__188__I5270 (.Y(N16693), .A(N16767), .B(N16789), .S0(N16800));
MXI2XL inst_cellmath__220__188__I5271 (.Y(N16727), .A(N16673), .B(N16662), .S0(N16800));
MXI2XL inst_cellmath__220__188__I5279 (.Y(N665), .A(N16798), .B(N16680), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5280 (.Y(N666), .A(N16708), .B(N16752), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5281 (.Y(N667), .A(N16780), .B(N16820), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5282 (.Y(N668), .A(N16689), .B(N16731), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5283 (.Y(N669), .A(N16761), .B(N16798), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5284 (.Y(N670), .A(N16666), .B(N16708), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5285 (.Y(N671), .A(N16739), .B(N16780), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5286 (.Y(N672), .A(N16808), .B(N16689), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5287 (.Y(N673), .A(N16717), .B(N16761), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5288 (.Y(N674), .A(N16788), .B(N16666), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5289 (.Y(N675), .A(N16699), .B(N16739), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5291 (.Y(N677), .A(N16676), .B(N16717), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5292 (.Y(N678), .A(N16711), .B(N16788), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5293 (.Y(N679), .A(N16750), .B(N16699), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5294 (.Y(N680), .A(N16783), .B(N16770), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5295 (.Y(N681), .A(N16817), .B(N16676), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5296 (.Y(N682), .A(N16693), .B(N16711), .S0(N16725));
MXI2XL inst_cellmath__220__188__I5297 (.Y(N683), .A(N16727), .B(N16750), .S0(N16725));
OR2XL cynw_cm_float_cos_I5304 (.Y(N709), .A(N16991), .B(N16722));
OR2XL cynw_cm_float_cos_I5305 (.Y(N710), .A(N16991), .B(N16759));
OR2XL cynw_cm_float_cos_I5306 (.Y(N711), .A(N16991), .B(inst_cellmath__215[2]));
OR2XL cynw_cm_float_cos_I5307 (.Y(N712), .A(N16991), .B(inst_cellmath__215[3]));
OR2XL cynw_cm_float_cos_I5308 (.Y(N713), .A(N16991), .B(inst_cellmath__215[4]));
NOR2XL inst_cellmath__223__199__I5357 (.Y(N17141), .A(inst_cellmath__42[6]), .B(inst_cellmath__19));
NOR4BBX1 inst_cellmath__223__199__I10822 (.Y(x[31]), .AN(N17141), .BN(N493), .C(inst_cellmath__42[8]), .D(inst_cellmath__42[7]));
OR2XL cynw_cm_float_cos_I5361 (.Y(N585), .A(inst_cellmath__68), .B(N16343));
NAND2BXL cynw_cm_float_cos_I5362 (.Y(N595), .AN(inst_cellmath__19), .B(N585));
NAND2XL cynw_cm_float_cos_I5364 (.Y(N594), .A(N17163), .B(inst_cellmath__68));
INVXL inst_cellmath__228_0_I5365 (.Y(N17178), .A(N741));
AO22XL inst_cellmath__228_0_I5366 (.Y(x[23]), .A0(N741), .A1(N594), .B0(N17178), .B1(N709));
AO22XL inst_cellmath__228_0_I5367 (.Y(x[24]), .A0(N741), .A1(N594), .B0(N17178), .B1(N710));
AO22XL inst_cellmath__228_0_I5368 (.Y(x[25]), .A0(N741), .A1(N594), .B0(N17178), .B1(N711));
AO22XL inst_cellmath__228_0_I5369 (.Y(x[26]), .A0(N741), .A1(N594), .B0(N17178), .B1(N712));
AO22XL inst_cellmath__228_0_I5370 (.Y(x[27]), .A0(N741), .A1(N594), .B0(N17178), .B1(N713));
OR2XL inst_cellmath__228_0_I5371 (.Y(x[28]), .A(N594), .B(N17178));
AND2XL inst_cellmath__228_0_I5373 (.Y(x[30]), .A(N595), .B(N741));
OR3XL inst_cellmath__231_0_I10823 (.Y(N17239), .A(N16991), .B(N16725), .C(N16680));
OR3XL inst_cellmath__231_0_I10557 (.Y(N17256), .A(N16991), .B(N16725), .C(N16752));
OR3XL inst_cellmath__231_0_I10537 (.Y(N17198), .A(N16991), .B(N16725), .C(N16820));
OR3XL inst_cellmath__231_0_I10550 (.Y(N17213), .A(N16991), .B(N16725), .C(N16731));
NAND2BXL inst_cellmath__231_0_I10482 (.Y(N17230), .AN(N16991), .B(N665));
NAND2BXL inst_cellmath__231_0_I10543 (.Y(N17247), .AN(N16991), .B(N666));
NAND2BXL inst_cellmath__231_0_I10476 (.Y(N17263), .AN(N16991), .B(N667));
NAND2BXL inst_cellmath__231_0_I10524 (.Y(N17205), .AN(N16991), .B(N668));
NAND2BXL inst_cellmath__231_0_I10458 (.Y(N17220), .AN(N16991), .B(N669));
NAND2BXL inst_cellmath__231_0_I10470 (.Y(N17237), .AN(N16991), .B(N670));
NAND2BXL inst_cellmath__231_0_I10500 (.Y(N17254), .AN(N16991), .B(N671));
NAND2BXL inst_cellmath__231_0_I10530 (.Y(N17270), .AN(N16991), .B(N672));
NAND2BXL inst_cellmath__231_0_I10506 (.Y(N17211), .AN(N16991), .B(N673));
NAND2BXL inst_cellmath__231_0_I10494 (.Y(N17227), .AN(N16991), .B(N674));
NAND2BXL inst_cellmath__231_0_I10512 (.Y(N17244), .AN(N16991), .B(N675));
NAND2BXL inst_cellmath__231_0_I10440 (.Y(N17202), .AN(N16991), .B(N677));
NAND2BXL inst_cellmath__231_0_I10434 (.Y(N17217), .AN(N16991), .B(N678));
NAND2BXL inst_cellmath__231_0_I10464 (.Y(N17234), .AN(N16991), .B(N679));
NAND2BXL inst_cellmath__231_0_I10488 (.Y(N17251), .AN(N16991), .B(N680));
NAND2BXL inst_cellmath__231_0_I10452 (.Y(N17267), .AN(N16991), .B(N681));
NAND2BXL inst_cellmath__231_0_I10428 (.Y(N17207), .AN(N16991), .B(N682));
NAND2BXL inst_cellmath__231_0_I10446 (.Y(N17223), .AN(N16991), .B(N683));
MXI2XL inst_cellmath__231_0_I5398 (.Y(x[0]), .A(N17239), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5399 (.Y(x[1]), .A(N17256), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5400 (.Y(x[2]), .A(N17198), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5401 (.Y(x[3]), .A(N17213), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5402 (.Y(x[4]), .A(N17230), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5403 (.Y(x[5]), .A(N17247), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5404 (.Y(x[6]), .A(N17263), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5405 (.Y(x[7]), .A(N17205), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5406 (.Y(x[8]), .A(N17220), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5407 (.Y(x[9]), .A(N17237), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5408 (.Y(x[10]), .A(N17254), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5409 (.Y(x[11]), .A(N17270), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5410 (.Y(x[12]), .A(N17211), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5411 (.Y(x[13]), .A(N17227), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5412 (.Y(x[14]), .A(N17244), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5414 (.Y(x[16]), .A(N17202), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5415 (.Y(x[17]), .A(N17217), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5416 (.Y(x[18]), .A(N17234), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5417 (.Y(x[19]), .A(N17251), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5418 (.Y(x[20]), .A(N17267), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5419 (.Y(x[21]), .A(N17207), .B(N17163), .S0(N741));
MXI2XL inst_cellmath__231_0_I5420 (.Y(x[22]), .A(N17223), .B(N17163), .S0(N741));
assign inst_cellmath__42[0] = 1'B0;
assign inst_cellmath__42[2] = 1'B0;
assign inst_cellmath__42[4] = 1'B0;
assign inst_cellmath__195[2] = 1'B0;
assign inst_cellmath__195[3] = 1'B0;
assign inst_cellmath__195[4] = 1'B0;
assign inst_cellmath__195[5] = 1'B0;
assign inst_cellmath__197[0] = 1'B0;
assign inst_cellmath__197[2] = 1'B0;
assign inst_cellmath__197[4] = 1'B0;
assign inst_cellmath__197[7] = 1'B0;
assign inst_cellmath__197[8] = 1'B0;
assign inst_cellmath__197[9] = 1'B0;
assign inst_cellmath__197[10] = 1'B0;
assign inst_cellmath__197[11] = 1'B0;
assign inst_cellmath__197[12] = 1'B0;
assign inst_cellmath__197[13] = 1'B0;
assign inst_cellmath__197[14] = 1'B0;
assign inst_cellmath__197[15] = 1'B0;
assign inst_cellmath__197[17] = 1'B0;
assign inst_cellmath__197[18] = 1'B0;
assign inst_cellmath__197[19] = 1'B0;
assign inst_cellmath__197[20] = 1'B1;
assign inst_cellmath__198[0] = 1'B0;
assign inst_cellmath__198[1] = 1'B0;
assign inst_cellmath__198[2] = 1'B0;
assign inst_cellmath__198[3] = 1'B0;
assign inst_cellmath__198[4] = 1'B0;
assign inst_cellmath__198[5] = 1'B0;
assign inst_cellmath__198[6] = 1'B0;
assign inst_cellmath__198[7] = 1'B0;
assign inst_cellmath__198[8] = 1'B0;
assign inst_cellmath__198[9] = 1'B0;
assign inst_cellmath__198[10] = 1'B0;
assign inst_cellmath__198[11] = 1'B0;
assign inst_cellmath__198[12] = 1'B0;
assign inst_cellmath__198[13] = 1'B0;
assign inst_cellmath__198[14] = 1'B0;
assign inst_cellmath__198[15] = 1'B0;
assign inst_cellmath__198[16] = 1'B0;
assign inst_cellmath__198[17] = 1'B0;
assign inst_cellmath__201[0] = 1'B0;
assign inst_cellmath__201[1] = 1'B0;
assign inst_cellmath__201[2] = 1'B0;
assign inst_cellmath__201[3] = 1'B0;
assign inst_cellmath__201[4] = 1'B0;
assign inst_cellmath__201[5] = 1'B0;
assign inst_cellmath__201[6] = 1'B0;
assign inst_cellmath__201[7] = 1'B0;
assign inst_cellmath__201[8] = 1'B0;
assign inst_cellmath__201[9] = 1'B0;
assign inst_cellmath__201[10] = 1'B0;
assign inst_cellmath__201[11] = 1'B0;
assign inst_cellmath__201[12] = 1'B0;
assign inst_cellmath__201[13] = 1'B0;
assign inst_cellmath__201[14] = 1'B0;
assign inst_cellmath__201[15] = 1'B0;
assign inst_cellmath__201[16] = 1'B0;
assign inst_cellmath__201[17] = 1'B0;
assign inst_cellmath__201[18] = 1'B0;
assign inst_cellmath__201[19] = 1'B0;
assign inst_cellmath__201[20] = 1'B0;
assign inst_cellmath__201[21] = 1'B0;
assign inst_cellmath__201[22] = 1'B0;
assign inst_cellmath__201[23] = 1'B0;
assign inst_cellmath__201[24] = 1'B0;
assign inst_cellmath__201[48] = 1'B0;
assign inst_cellmath__203__W0[0] = 1'B0;
assign inst_cellmath__203__W0[20] = 1'B0;
assign inst_cellmath__203__W0[21] = 1'B0;
assign inst_cellmath__203__W0[22] = 1'B0;
assign inst_cellmath__203__W0[23] = 1'B0;
assign inst_cellmath__203__W0[43] = 1'B1;
assign inst_cellmath__203__W0[44] = 1'B1;
assign inst_cellmath__203__W0[45] = 1'B1;
assign inst_cellmath__203__W0[46] = 1'B1;
assign inst_cellmath__203__W1[0] = 1'B0;
assign inst_cellmath__203__W1[20] = 1'B0;
assign inst_cellmath__203__W1[21] = 1'B0;
assign inst_cellmath__203__W1[22] = 1'B0;
assign inst_cellmath__203__W1[23] = 1'B0;
assign inst_cellmath__203__W1[43] = 1'B0;
assign inst_cellmath__203__W1[44] = 1'B0;
assign inst_cellmath__203__W1[45] = 1'B0;
assign inst_cellmath__203__W1[46] = 1'B0;
assign inst_cellmath__210[23] = 1'B0;
assign inst_cellmath__210[24] = 1'B0;
assign inst_cellmath__210[25] = 1'B0;
assign inst_cellmath__210[26] = 1'B0;
assign inst_cellmath__210[27] = 1'B0;
assign inst_cellmath__210[28] = 1'B0;
assign inst_cellmath__210[29] = 1'B0;
assign inst_cellmath__210[30] = 1'B0;
assign inst_cellmath__215[1] = 1'B0;
assign x[29] = x[28];
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  v7jzSg/arBs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



