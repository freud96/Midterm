/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 11:19:26 CST (+0800), Sunday 24 April 2022
    Configured on: ws45
    Configured by: m110061422 (m110061422)
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadtool/cadence/STRATUS/cur/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadtool/cadence/STRATUS/STRATUS_19.12.100/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module DFT_compute_cynw_cm_float_mul_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
output [31:0] x;
wire  inst_cellmath__17,
	inst_cellmath__18,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23,
	inst_cellmath__24,
	inst_cellmath__25,
	inst_cellmath__26,
	inst_cellmath__29,
	inst_cellmath__33;
wire [9:0] inst_cellmath__34;
wire  inst_cellmath__41,
	inst_cellmath__42;
wire [47:0] inst_cellmath__43;
wire [7:0] inst_cellmath__50;
wire N269,N270,N272,N273,N274,N1736,N1740 
	,N1758,N1762,N1779,N1787,N1793,N1795,N1798,N1800 
	,N1808,N1810,N1814,N1820,N1859,N1863,N1881,N1885 
	,N1902,N1904,N1906,N1910,N1916,N1921,N1933,N1937 
	,N1941,N1943,N1999,N2011,N2012,N2013,N2014,N2015 
	,N2016,N2018,N2019,N2020,N2021,N2022,N2023,N2024 
	,N2026,N2027,N2028,N2029,N2030,N2032,N2034,N2036 
	,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2045 
	,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053 
	,N2055,N2056,N2057,N2059,N2060,N2061,N2063,N2064 
	,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072 
	,N2073,N2075,N2076,N2077,N2079,N2080,N2081,N2082 
	,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090 
	,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098 
	,N2099,N2101,N2102,N2103,N2104,N2105,N2106,N2107 
	,N2108,N2109,N2110,N2111,N2113,N2114,N2115,N2116 
	,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124 
	,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132 
	,N2133,N2134,N2135,N2136,N2138,N2139,N2140,N2141 
	,N2142,N2143,N2144,N2145,N2146,N2147,N2149,N2151 
	,N2152,N2153,N2154,N2156,N2157,N2158,N2159,N2160 
	,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168 
	,N2169,N2171,N2172,N2173,N2174,N2175,N2176,N2178 
	,N2179,N2181,N2182,N2183,N2184,N2185,N2186,N2187 
	,N2188,N2189,N2190,N2191,N2193,N2194,N2195,N2196 
	,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204 
	,N2205,N2206,N2208,N2209,N2210,N2211,N2212,N2213 
	,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2222 
	,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230 
	,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238 
	,N2239,N2240,N2241,N2244,N2245,N2246,N2247,N2248 
	,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256 
	,N2257,N2258,N2259,N2260,N2263,N2264,N2265,N2266 
	,N2267,N2268,N2269,N2270,N2272,N2273,N2274,N2275 
	,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283 
	,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291 
	,N2292,N2293,N2294,N2295,N2296,N2297,N2299,N2300 
	,N2301,N2302,N2303,N2304,N2305,N2306,N2308,N2309 
	,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317 
	,N2318,N2319,N2321,N2322,N2323,N2324,N2325,N2326 
	,N2327,N2329,N2330,N2331,N2332,N2333,N2334,N2335 
	,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344 
	,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352 
	,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360 
	,N2361,N2362,N2363,N2365,N2366,N2367,N2368,N2369 
	,N2370,N2371,N2372,N2373,N2374,N2375,N2377,N2379 
	,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387 
	,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395 
	,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403 
	,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411 
	,N2412,N2415,N2416,N2417,N2418,N2419,N2420,N2421 
	,N2422,N2423,N2424,N2426,N2427,N2428,N2429,N2430 
	,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438 
	,N2440,N2441,N2443,N2444,N2445,N2447,N2448,N2449 
	,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2459 
	,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467 
	,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475 
	,N2476,N2477,N2478,N2479,N2480,N2482,N2483,N2484 
	,N2485,N2486,N2487,N2488,N2490,N2491,N2492,N2493 
	,N2494,N2495,N2496,N2497,N2499,N2500,N2501,N2502 
	,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510 
	,N2511,N2512,N2514,N2515,N2516,N2517,N2518,N2520 
	,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528 
	,N2530,N2531,N2532,N2534,N2535,N2536,N2537,N2538 
	,N2539,N2540,N2541,N2543,N2544,N2545,N2546,N2547 
	,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555 
	,N2556,N2558,N2559,N2560,N2561,N2562,N2563,N2564 
	,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573 
	,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2582 
	,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2591 
	,N2593,N2596,N2597,N2598,N2599,N2602,N2604,N2605 
	,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613 
	,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621 
	,N2622,N2623,N2625,N2626,N2627,N2628,N2629,N2630 
	,N2631,N2632,N2633,N2634,N2636,N2637,N2638,N2639 
	,N2640,N2641,N2642,N2644,N2645,N2646,N2647,N2648 
	,N2649,N2650,N2652,N2653,N2654,N2655,N2656,N2657 
	,N2658,N2660,N2661,N2662,N2663,N2664,N2665,N2666 
	,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674 
	,N2675,N2677,N2678,N2680,N2681,N2682,N2683,N2684 
	,N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692 
	,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2701 
	,N2703,N2704,N2705,N2706,N2707,N2709,N2710,N2711 
	,N2712,N2713,N2714,N2715,N2717,N2719,N2720,N2721 
	,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729 
	,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737 
	,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745 
	,N2746,N2747,N2748,N2749,N2750,N2751,N2753,N2754 
	,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762 
	,N2763,N2764,N2765,N2766,N2767,N2768,N2770,N2771 
	,N2772,N2774,N2775,N2777,N2778,N2779,N2780,N2781 
	,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789 
	,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2798 
	,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2807 
	,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815 
	,N2816,N2818,N2819,N2820,N2821,N2822,N2823,N2824 
	,N2825,N2826,N2827,N2828,N2829,N2831,N2832,N2833 
	,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841 
	,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849 
	,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857 
	,N2858,N2860,N2862,N2863,N2865,N2866,N2867,N2871 
	,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879 
	,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887 
	,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895 
	,N2896,N2897,N2898,N2899,N2901,N2902,N2903,N2904 
	,N2905,N2906,N2907,N2908,N2909,N2910,N2912,N2913 
	,N2914,N2915,N2916,N2918,N2919,N2920,N2922,N2923 
	,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2932 
	,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940 
	,N2941,N2942,N2943,N2944,N2945,N2946,N2948,N2949 
	,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957 
	,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2966 
	,N2967,N2968,N2969,N2970,N2971,N2973,N2974,N2975 
	,N2978,N2979,N2980,N2982,N2983,N2984,N2985,N2986 
	,N2987,N2988,N2991,N2992,N2993,N2994,N2995,N2996 
	,N2997,N2998,N3000,N3001,N3002,N3003,N3004,N3005 
	,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3014 
	,N3015,N3016,N3018,N3019,N3020,N3021,N3022,N3023 
	,N3025,N3027,N3028,N3029,N3030,N3031,N3032,N3033 
	,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041 
	,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3050 
	,N3052,N3054,N3055,N3056,N3057,N3058,N3059,N3060 
	,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070 
	,N3071,N3073,N3074,N3075,N3076,N3077,N3078,N3079 
	,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087 
	,N3088,N3090,N3091,N3092,N3093,N3094,N3096,N3097 
	,N3098,N3099,N3101,N3102,N3103,N3104,N3106,N3107 
	,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115 
	,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123 
	,N3124,N3125,N3127,N3128,N3129,N3130,N3131,N3132 
	,N3133,N3134,N3136,N3139,N3140,N3141,N3142,N3143 
	,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151 
	,N3152,N3154,N3155,N3156,N3157,N3158,N3159,N3160 
	,N3161,N3162,N3164,N3165,N3166,N3167,N3168,N3169 
	,N3171,N3172,N3173,N3174,N3176,N3177,N3178,N3179 
	,N3180,N3181,N3182,N3183,N3185,N3186,N3187,N3188 
	,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196 
	,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204 
	,N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212 
	,N3213,N3214,N3215,N3216,N3218,N3219,N3220,N3221 
	,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229 
	,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237 
	,N3238,N3240,N3241,N3244,N3245,N3246,N3249,N3250 
	,N3251,N3252,N3253,N3254,N3255,N3256,N3258,N3259 
	,N3260,N3261,N3262,N3263,N3264,N3266,N3267,N3268 
	,N3269,N3270,N3271,N3273,N3274,N3275,N3276,N3277 
	,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285 
	,N3286,N3287,N3288,N3289,N3291,N3292,N3293,N3294 
	,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302 
	,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310 
	,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3319 
	,N3320,N3321,N3322,N3323,N3324,N3326,N3327,N3328 
	,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337 
	,N3338,N3339,N3340,N3341,N3342,N3343,N3344,N3345 
	,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353 
	,N3354,N3355,N3356,N3357,N3359,N3360,N3361,N3363 
	,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3372 
	,N3373,N3374,N3375,N3377,N3379,N3380,N3381,N3382 
	,N3383,N3384,N3385,N3386,N3387,N3388,N3390,N3391 
	,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399 
	,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407 
	,N3409,N3411,N3412,N3413,N3414,N3415,N3416,N3417 
	,N3418,N3419,N3420,N3422,N3423,N3425,N3426,N3427 
	,N3428,N3429,N3430,N3431,N3432,N3433,N3435,N3436 
	,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444 
	,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452 
	,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460 
	,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468 
	,N3469,N3470,N3471,N3472,N3473,N3475,N3476,N3477 
	,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485 
	,N3486,N3487,N3489,N3490,N3491,N3492,N3493,N3494 
	,N3495,N3497,N3498,N3499,N3500,N3501,N3502,N3503 
	,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511 
	,N3512,N3513,N3514,N3516,N3517,N3518,N3519,N3520 
	,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530 
	,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538 
	,N3539,N3542,N3543,N3544,N3545,N3546,N3547,N3548 
	,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556 
	,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564 
	,N3565,N3566,N3567,N3569,N3570,N3571,N3572,N3573 
	,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581 
	,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589 
	,N3590,N3591,N3592,N3593,N3594,N3596,N3597,N3598 
	,N3599,N3600,N3601,N3602,N3604,N3605,N3606,N3607 
	,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615 
	,N3616,N3618,N3619,N3620,N3621,N3623,N3624,N3626 
	,N3627,N3628,N3629,N3630,N3631,N3633,N3634,N3635 
	,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643 
	,N3644,N3646,N3647,N3648,N3649,N3650,N3651,N3652 
	,N3653,N3654,N3655,N3656,N3657,N3659,N3660,N3661 
	,N3662,N3663,N3664,N3666,N3667,N3668,N3669,N3670 
	,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678 
	,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687 
	,N3688,N3689,N3690,N3691,N3692,N3693,N3695,N3696 
	,N3697,N3698,N3699,N3700,N3701,N3702,N3705,N3706 
	,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714 
	,N3715,N3716,N3717,N3719,N3720,N3721,N3722,N3723 
	,N3724,N3725,N3726,N3727,N3728,N3729,N3730,N3731 
	,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3740 
	,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3749 
	,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757 
	,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765 
	,N3766,N3767,N3768,N3769,N3770,N3771,N3773,N3774 
	,N3775,N3776,N3777,N3778,N3779,N3781,N3784,N3785 
	,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793 
	,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802 
	,N3803,N3804,N3805,N3807,N3808,N3809,N3810,N3811 
	,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820 
	,N3821,N3822,N3823,N3824,N3826,N3827,N3828,N3829 
	,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837 
	,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845 
	,N3846,N3847,N3848,N3849,N3851,N3852,N3853,N3854 
	,N3855,N3856,N3857,N3858,N3861,N3862,N3863,N3864 
	,N3865,N3866,N3867,N3868,N3869,N3871,N3872,N3873 
	,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881 
	,N3882,N3883,N3885,N3887,N3888,N3889,N3890,N3892 
	,N3893,N3894,N3895,N3896,N3897,N3898,N3900,N3902 
	,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910 
	,N3911,N3912,N3913,N3914,N3915,N3916,N3917,N3918 
	,N3919,N3920,N3921,N3922,N3923,N3925,N3926,N3927 
	,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935 
	,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944 
	,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952 
	,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3961 
	,N3962,N3963,N3965,N3966,N3967,N3968,N3969,N3972 
	,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981 
	,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989 
	,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997 
	,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005 
	,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013 
	,N4014,N4016,N4017,N4018,N4019,N4020,N4021,N4022 
	,N4024,N4025,N4026,N4028,N4029,N4030,N4031,N4032 
	,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040 
	,N4041,N4042,N4043,N4045,N4046,N4047,N4048,N4051 
	,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060 
	,N4061,N4063,N4064,N4065,N4066,N4067,N4068,N4069 
	,N4070,N4071,N4072,N4074,N4075,N4076,N4078,N4079 
	,N4080,N4081,N4082,N4083,N4084,N4085,N4087,N4088 
	,N4089,N4090,N4091,N4092,N4093,N4094,N4096,N4097 
	,N4098,N4099,N4100,N4101,N4102,N4103,N4104,N4105 
	,N6156,N6163,N6169,N6175,N6176,N6177,N6178,N6180 
	,N6181,N6183,N6184,N6186,N6188,N6189,N6190,N6192 
	,N6193,N6196,N6197,N6198,N6199,N6200,N6201,N6202 
	,N6203,N6204,N6206,N6207,N6210,N6211,N6213,N6215 
	,N6218,N6220,N6222,N6223,N6224,N6226,N6227,N6229 
	,N6230,N6231,N6232,N6233,N6234,N6236,N6237,N6240 
	,N6242,N6244,N6245,N6247,N6248,N6249,N6251,N6252 
	,N6253,N6254,N6256,N6257,N6258,N6259,N6261,N6263 
	,N6337,N6342,N6349,N6355,N6367,N6374,N6381,N6386 
	,N6389,N6417,N6424,N6426,N6437,N6439,N6457,N6469 
	,N6480,N6494,N6503,N6504,N6505,N6508,N6513,N6524 
	,N6525,N6551,N6564,N6567,N6571,N6575,N6578,N6581 
	,N6583,N6584,N6588,N6593,N6596,N6600,N6604,N6608 
	,N6610,N6613,N6618,N6625,N6629,N6633,N6635,N6636 
	,N6639,N6640,N6647,N6652,N6654,N6659,N6663,N6666 
	,N6669,N6670,N6675,N6680,N6683,N6687,N9354,N9370 
	,N9371,N9378,N9379,N9380,N9381,N9391,N9399,N9406 
	,N9410,N9417,N9426,N18785,N18795,N18799,N18814,N18818 
	,N18820,N18823,N18825,N18827,N18836,N18839,N18841,N18846 
	,N18848,N18857,N18860,N18886,N18898,N18901,N18904,N18917 
	,N18923;
XNOR2X1 cynw_cm_float_mul_I4111 (.Y(inst_cellmath__33), .A(a_sign), .B(b_sign));
OR4X1 inst_cellmath__26__8__I11214 (.Y(N1736), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__26__8__I11215 (.Y(N1740), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL inst_cellmath__26__8__I293 (.Y(inst_cellmath__26), .A(N1736), .B(N1740));
AND4XL inst_cellmath__17_0_I11216 (.Y(N1758), .A(a_exp[0]), .B(a_exp[1]), .C(a_exp[7]), .D(a_exp[6]));
AND4XL inst_cellmath__17_0_I11217 (.Y(N1762), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND2XL inst_cellmath__17_0_I300 (.Y(inst_cellmath__17), .A(N1758), .B(N1762));
NOR2XL inst_cellmath__19__5__I301 (.Y(N1808), .A(a_man[0]), .B(a_man[1]));
NOR2XL inst_cellmath__19__5__I309 (.Y(N1795), .A(a_man[8]), .B(a_man[7]));
CLKINVX8 inst_cellmath__19__5__I312 (.Y(N1779), .A(a_man[2]));
OR4X1 inst_cellmath__19__5__I11218 (.Y(N1800), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__19__5__I11219 (.Y(N1810), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__19__5__I11220 (.Y(N1820), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
OR4X1 inst_cellmath__19__5__I11222 (.Y(N1793), .A(a_man[6]), .B(a_man[4]), .C(a_man[5]), .D(a_man[3]));
NOR4BX1 inst_cellmath__19__5__I11223 (.Y(N1798), .AN(N1795), .B(a_man[10]), .C(N1793), .D(a_man[9]));
NOR2XL inst_cellmath__19__5__I320 (.Y(N1814), .A(N1810), .B(N1820));
NAND3XL hyperpropagate_4_1_A_I4228 (.Y(N9391), .A(N1779), .B(N1808), .C(N1814));
NOR2XL hyperpropagate_4_1_A_I4229 (.Y(N1787), .A(N1800), .B(N9391));
NAND2XL inst_cellmath__19__5__I323 (.Y(inst_cellmath__19), .A(N1798), .B(N1787));
NOR2XL cynw_cm_float_mul_I324 (.Y(inst_cellmath__23), .A(inst_cellmath__17), .B(inst_cellmath__19));
OR4X1 inst_cellmath__25__7__I11224 (.Y(N1859), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__25__7__I11225 (.Y(N1863), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__25__7__I333 (.Y(inst_cellmath__25), .A(N1859), .B(N1863));
AND4XL inst_cellmath__18_0_I11226 (.Y(N1881), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[7]), .D(b_exp[6]));
AND4XL inst_cellmath__18_0_I11227 (.Y(N1885), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND2XL inst_cellmath__18_0_I340 (.Y(inst_cellmath__18), .A(N1881), .B(N1885));
NOR2XL inst_cellmath__20__6__I342 (.Y(N1941), .A(b_man[22]), .B(b_man[21]));
NOR2XL inst_cellmath__20__6__I343 (.Y(N1904), .A(b_man[20]), .B(b_man[19]));
CLKINVX8 inst_cellmath__20__6__I352 (.Y(N1902), .A(b_man[2]));
CLKINVX6 inst_cellmath__20__6__I4086 (.Y(N9370), .A(N1902));
CLKINVX8 inst_cellmath__20__6__I4087 (.Y(N9371), .A(N9370));
OR4X1 inst_cellmath__20__6__I11229 (.Y(N1933), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__20__6__I11230 (.Y(N1943), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR2XL inst_cellmath__20__6__I360 (.Y(N1937), .A(N1933), .B(N1943));
NAND3XL hyperpropagate_4_1_A_I4230 (.Y(N9399), .A(N1941), .B(N1904), .C(N1937));
NOR4BX1 hyperpropagate_4_1_A_I11233 (.Y(N1910), .AN(N9371), .B(b_man[0]), .C(N9399), .D(b_man[1]));
OR4X1 inst_cellmath__20__6__I11231 (.Y(N1906), .A(b_man[10]), .B(b_man[8]), .C(b_man[9]), .D(b_man[7]));
OR4X1 inst_cellmath__20__6__I11232 (.Y(N1916), .A(b_man[6]), .B(b_man[4]), .C(b_man[5]), .D(b_man[3]));
NOR2XL inst_cellmath__20__6__I362 (.Y(N1921), .A(N1906), .B(N1916));
NAND2XL inst_cellmath__20__6__I363 (.Y(inst_cellmath__20), .A(N1921), .B(N1910));
NOR2XL cynw_cm_float_mul_I364 (.Y(inst_cellmath__24), .A(inst_cellmath__18), .B(inst_cellmath__20));
NOR2BX1 cynw_cm_float_mul_I4115 (.Y(inst_cellmath__21), .AN(inst_cellmath__19), .B(inst_cellmath__17));
NOR2BX1 cynw_cm_float_mul_I4116 (.Y(inst_cellmath__22), .AN(inst_cellmath__20), .B(inst_cellmath__18));
AOI211XL inst_cellmath__29_0_I4169 (.Y(N1999), .A0(inst_cellmath__26), .A1(inst_cellmath__23), .B0(inst_cellmath__21), .C0(inst_cellmath__22));
OAI2BB1X1 inst_cellmath__29_0_I4118 (.Y(inst_cellmath__29), .A0N(inst_cellmath__25), .A1N(inst_cellmath__24), .B0(N1999));
NOR2XL cynw_cm_float_mul_I377 (.Y(x[31]), .A(inst_cellmath__33), .B(inst_cellmath__29));
CLKINVX4 inst_cellmath__43_0_I378 (.Y(N3614), .A(b_man[0]));
CLKINVX6 inst_cellmath__43_0_I380 (.Y(N3075), .A(b_man[1]));
CLKINVX4 inst_cellmath__43_0_I384 (.Y(N4097), .A(b_man[3]));
CLKINVX6 inst_cellmath__43_0_I385 (.Y(N3571), .A(b_man[4]));
CLKINVX6 inst_cellmath__43_0_I386 (.Y(N3029), .A(b_man[5]));
CLKINVX6 inst_cellmath__43_0_I387 (.Y(N2490), .A(b_man[6]));
CLKINVX8 inst_cellmath__43_0_I388 (.Y(N4055), .A(b_man[7]));
CLKINVX12 inst_cellmath__43_0_I390 (.Y(N3526), .A(b_man[8]));
CLKINVX8 inst_cellmath__43_0_I392 (.Y(N2984), .A(b_man[9]));
CLKINVX8 inst_cellmath__43_0_I394 (.Y(N2451), .A(b_man[10]));
CLKINVX12 inst_cellmath__43_0_I396 (.Y(N4008), .A(b_man[11]));
CLKINVX12 inst_cellmath__43_0_I398 (.Y(N3479), .A(b_man[12]));
CLKINVX8 inst_cellmath__43_0_I401 (.Y(N2940), .A(b_man[13]));
CLKINVX20 inst_cellmath__43_0_I403 (.Y(N2405), .A(b_man[14]));
CLKINVX12 inst_cellmath__43_0_I405 (.Y(N3963), .A(b_man[15]));
CLKINVX12 inst_cellmath__43_0_I407 (.Y(N3437), .A(b_man[16]));
CLKINVX12 inst_cellmath__43_0_I408 (.Y(N2895), .A(b_man[17]));
CLKINVX6 inst_cellmath__43_0_I410 (.Y(N2360), .A(b_man[18]));
CLKINVX8 inst_cellmath__43_0_I411 (.Y(N3920), .A(b_man[19]));
CLKINVX8 inst_cellmath__43_0_I412 (.Y(N3391), .A(b_man[20]));
CLKINVX6 inst_cellmath__43_0_I413 (.Y(N2849), .A(b_man[21]));
CLKINVX6 inst_cellmath__43_0_I414 (.Y(N2317), .A(b_man[22]));
CLKINVX8 inst_cellmath__43_0_I415 (.Y(N3878), .A(a_man[0]));
NOR2XL inst_cellmath__43_0_I419 (.Y(N4036), .A(N3878), .B(N9371));
NOR2XL inst_cellmath__43_0_I420 (.Y(N2855), .A(N3878), .B(N4097));
NOR2XL inst_cellmath__43_0_I421 (.Y(N3769), .A(N3878), .B(N3571));
NOR2XL inst_cellmath__43_0_I422 (.Y(N2589), .A(N3878), .B(N3029));
NOR2XL inst_cellmath__43_0_I423 (.Y(N3511), .A(N3878), .B(N2490));
NOR2XL inst_cellmath__43_0_I424 (.Y(N2323), .A(N3878), .B(N4055));
NOR2XL inst_cellmath__43_0_I425 (.Y(N3236), .A(N3878), .B(N3526));
NOR2XL inst_cellmath__43_0_I426 (.Y(N2059), .A(N3878), .B(N2984));
NOR2XL inst_cellmath__43_0_I427 (.Y(N2966), .A(N3878), .B(N2451));
NOR2XL inst_cellmath__43_0_I428 (.Y(N3881), .A(N3878), .B(N4008));
NOR2XL inst_cellmath__43_0_I429 (.Y(N2698), .A(N3878), .B(N3479));
NOR2XL inst_cellmath__43_0_I430 (.Y(N3627), .A(N3878), .B(N2940));
NOR2XL inst_cellmath__43_0_I431 (.Y(N2435), .A(N3878), .B(N2405));
NOR2XL inst_cellmath__43_0_I432 (.Y(N3351), .A(N3878), .B(N3963));
NOR2XL inst_cellmath__43_0_I433 (.Y(N2171), .A(N3878), .B(N3437));
NOR2XL inst_cellmath__43_0_I434 (.Y(N3086), .A(N3878), .B(N2895));
NOR2XL inst_cellmath__43_0_I435 (.Y(N3996), .A(N3878), .B(N2360));
NOR2XL inst_cellmath__43_0_I436 (.Y(N2811), .A(N3878), .B(N3920));
NOR2X2 inst_cellmath__43_0_I437 (.Y(N3731), .A(N3878), .B(N3391));
NOR2XL inst_cellmath__43_0_I438 (.Y(N2545), .A(N3878), .B(N2849));
NOR2X1 inst_cellmath__43_0_I439 (.Y(N3464), .A(N3878), .B(N2317));
INVXL inst_cellmath__43_0_I440 (.Y(N2279), .A(N3878));
CLKINVX8 inst_cellmath__43_0_I441 (.Y(N3347), .A(a_man[1]));
NOR2XL inst_cellmath__43_0_I444 (.Y(N2843), .A(N3347), .B(N3075));
NOR2XL inst_cellmath__43_0_I445 (.Y(N3760), .A(N3347), .B(N9371));
NOR2XL inst_cellmath__43_0_I446 (.Y(N2578), .A(N3347), .B(N4097));
NOR2XL inst_cellmath__43_0_I447 (.Y(N3501), .A(N3347), .B(N3571));
NOR2XL inst_cellmath__43_0_I448 (.Y(N2313), .A(N3347), .B(N3029));
NOR2XL inst_cellmath__43_0_I449 (.Y(N3229), .A(N3347), .B(N2490));
NOR2XL inst_cellmath__43_0_I450 (.Y(N2048), .A(N3347), .B(N4055));
NOR2XL inst_cellmath__43_0_I451 (.Y(N2959), .A(N3347), .B(N3526));
NOR2XL inst_cellmath__43_0_I452 (.Y(N3871), .A(N3347), .B(N2984));
NOR2XL inst_cellmath__43_0_I453 (.Y(N2689), .A(N3347), .B(N2451));
NOR2XL inst_cellmath__43_0_I454 (.Y(N3616), .A(N3347), .B(N4008));
NOR2XL inst_cellmath__43_0_I455 (.Y(N2426), .A(N3347), .B(N3479));
NOR2XL inst_cellmath__43_0_I456 (.Y(N3340), .A(N3347), .B(N2940));
NOR2XL inst_cellmath__43_0_I457 (.Y(N2163), .A(N3347), .B(N2405));
NOR2XL inst_cellmath__43_0_I458 (.Y(N3076), .A(N3347), .B(N3963));
NOR2XL inst_cellmath__43_0_I459 (.Y(N3986), .A(N3347), .B(N3437));
NOR2XL inst_cellmath__43_0_I460 (.Y(N2801), .A(N3347), .B(N2895));
NOR2XL inst_cellmath__43_0_I461 (.Y(N3722), .A(N3347), .B(N2360));
NOR2X2 inst_cellmath__43_0_I462 (.Y(N2534), .A(N3347), .B(N3920));
NOR2XL inst_cellmath__43_0_I463 (.Y(N3457), .A(N3347), .B(N3391));
NOR2XL inst_cellmath__43_0_I464 (.Y(N2266), .A(N3347), .B(N2849));
NOR2X1 inst_cellmath__43_0_I465 (.Y(N3187), .A(N3347), .B(N2317));
INVXL inst_cellmath__43_0_I466 (.Y(N4101), .A(N3347));
NOR2XL inst_cellmath__43_0_I469 (.Y(N3752), .A(N1779), .B(N3614));
NOR2XL inst_cellmath__43_0_I470 (.Y(N2570), .A(N1779), .B(N3075));
NOR2XL inst_cellmath__43_0_I471 (.Y(N3491), .A(N1779), .B(N9371));
NOR2XL inst_cellmath__43_0_I472 (.Y(N2302), .A(N1779), .B(N4097));
NOR2XL inst_cellmath__43_0_I473 (.Y(N3220), .A(N1779), .B(N3571));
NOR2XL inst_cellmath__43_0_I474 (.Y(N2038), .A(N1779), .B(N3029));
NOR2XL inst_cellmath__43_0_I475 (.Y(N2951), .A(N1779), .B(N2490));
NOR2XL inst_cellmath__43_0_I476 (.Y(N3863), .A(N1779), .B(N4055));
NOR2XL inst_cellmath__43_0_I477 (.Y(N2680), .A(N1779), .B(N3526));
NOR2XL inst_cellmath__43_0_I478 (.Y(N3606), .A(N1779), .B(N2984));
NOR2XL inst_cellmath__43_0_I479 (.Y(N2418), .A(N1779), .B(N2451));
NOR2XL inst_cellmath__43_0_I480 (.Y(N3332), .A(N1779), .B(N4008));
NOR2XL inst_cellmath__43_0_I481 (.Y(N2152), .A(N1779), .B(N3479));
NOR2XL inst_cellmath__43_0_I482 (.Y(N3066), .A(N1779), .B(N2940));
NOR2XL inst_cellmath__43_0_I483 (.Y(N3976), .A(N1779), .B(N2405));
NOR2XL inst_cellmath__43_0_I484 (.Y(N2791), .A(N1779), .B(N3963));
NOR2XL inst_cellmath__43_0_I485 (.Y(N3715), .A(N1779), .B(N3437));
NOR2XL inst_cellmath__43_0_I486 (.Y(N2524), .A(N2895), .B(N1779));
NOR2X1 inst_cellmath__43_0_I487 (.Y(N3449), .A(N1779), .B(N2360));
NOR2X1 inst_cellmath__43_0_I488 (.Y(N2256), .A(N3920), .B(N1779));
NOR2X2 inst_cellmath__43_0_I489 (.Y(N3176), .A(N3391), .B(N1779));
NOR2X1 inst_cellmath__43_0_I490 (.Y(N4090), .A(N1779), .B(N2849));
NOR2X1 inst_cellmath__43_0_I491 (.Y(N2906), .A(N2317), .B(N1779));
INVXL inst_cellmath__43_0_I492 (.Y(N3817), .A(N1779));
CLKINVX8 inst_cellmath__43_0_I493 (.Y(N2274), .A(a_man[3]));
NOR2XL inst_cellmath__43_0_I495 (.Y(N3480), .A(N2274), .B(N3614));
NOR2XL inst_cellmath__43_0_I496 (.Y(N2292), .A(N2274), .B(N3075));
NOR2XL inst_cellmath__43_0_I497 (.Y(N3211), .A(N2274), .B(N9371));
NOR2XL inst_cellmath__43_0_I498 (.Y(N2027), .A(N2274), .B(N4097));
NOR2XL inst_cellmath__43_0_I499 (.Y(N2941), .A(N2274), .B(N3571));
NOR2XL inst_cellmath__43_0_I500 (.Y(N3852), .A(N2274), .B(N3029));
NOR2XL inst_cellmath__43_0_I501 (.Y(N2671), .A(N2274), .B(N2490));
NOR2XL inst_cellmath__43_0_I502 (.Y(N3598), .A(N2274), .B(N4055));
NOR2XL inst_cellmath__43_0_I503 (.Y(N2408), .A(N2274), .B(N3526));
NOR2XL inst_cellmath__43_0_I504 (.Y(N3321), .A(N2274), .B(N2984));
NOR2XL inst_cellmath__43_0_I505 (.Y(N2140), .A(N2274), .B(N2451));
NOR2XL inst_cellmath__43_0_I506 (.Y(N3056), .A(N2274), .B(N4008));
NOR2XL inst_cellmath__43_0_I507 (.Y(N3965), .A(N2274), .B(N3479));
NOR2XL inst_cellmath__43_0_I508 (.Y(N2779), .A(N2274), .B(N2940));
NOR2XL inst_cellmath__43_0_I509 (.Y(N3706), .A(N2274), .B(N2405));
NOR2XL inst_cellmath__43_0_I510 (.Y(N2515), .A(N2274), .B(N3963));
NOR2XL inst_cellmath__43_0_I511 (.Y(N3438), .A(N2274), .B(N3437));
NOR2X1 inst_cellmath__43_0_I512 (.Y(N2247), .A(N2895), .B(N2274));
NOR2X1 inst_cellmath__43_0_I513 (.Y(N3167), .A(N2274), .B(N2360));
NOR2X2 inst_cellmath__43_0_I514 (.Y(N4079), .A(N2274), .B(N3920));
NOR2XL inst_cellmath__43_0_I515 (.Y(N2898), .A(N2274), .B(N3391));
NOR2X2 inst_cellmath__43_0_I516 (.Y(N3809), .A(N2274), .B(N2849));
NOR2XL inst_cellmath__43_0_I517 (.Y(N2631), .A(N2274), .B(N2317));
INVXL inst_cellmath__43_0_I518 (.Y(N3553), .A(N2274));
CLKINVX12 inst_cellmath__43_0_I519 (.Y(N3833), .A(a_man[4]));
INVX8 inst_cellmath__43_0_I4094 (.Y(N9378), .A(N3833));
INVX12 inst_cellmath__43_0_I4095 (.Y(N9379), .A(N9378));
NOR2XL inst_cellmath__43_0_I521 (.Y(N3203), .A(N9379), .B(N3614));
NOR2XL inst_cellmath__43_0_I522 (.Y(N2019), .A(N9379), .B(N3075));
NOR2XL inst_cellmath__43_0_I523 (.Y(N2932), .A(N9379), .B(N9371));
NOR2XL inst_cellmath__43_0_I524 (.Y(N3844), .A(N9379), .B(N4097));
NOR2XL inst_cellmath__43_0_I525 (.Y(N2661), .A(N9379), .B(N3571));
NOR2XL inst_cellmath__43_0_I526 (.Y(N3589), .A(N9379), .B(N3029));
NOR2XL inst_cellmath__43_0_I527 (.Y(N2398), .A(N9379), .B(N2490));
NOR2XL inst_cellmath__43_0_I528 (.Y(N3311), .A(N9379), .B(N4055));
NOR2XL inst_cellmath__43_0_I529 (.Y(N2129), .A(N9379), .B(N3526));
NOR2XL inst_cellmath__43_0_I530 (.Y(N3043), .A(N9379), .B(N2984));
NOR2XL inst_cellmath__43_0_I531 (.Y(N3952), .A(N9379), .B(N2451));
NOR2XL inst_cellmath__43_0_I532 (.Y(N2766), .A(N9379), .B(N4008));
NOR2XL inst_cellmath__43_0_I533 (.Y(N3695), .A(N9379), .B(N3479));
NOR2XL inst_cellmath__43_0_I534 (.Y(N2506), .A(N9379), .B(N2940));
NOR2XL inst_cellmath__43_0_I535 (.Y(N3427), .A(N9379), .B(N2405));
NOR2XL inst_cellmath__43_0_I536 (.Y(N2237), .A(N3963), .B(N9379));
NOR2X2 inst_cellmath__43_0_I537 (.Y(N3156), .A(N3437), .B(N9379));
NOR2X1 inst_cellmath__43_0_I538 (.Y(N4069), .A(N2895), .B(N9379));
NOR2XL inst_cellmath__43_0_I539 (.Y(N2888), .A(N3833), .B(N2360));
NOR2X1 inst_cellmath__43_0_I540 (.Y(N3800), .A(N3920), .B(N3833));
NOR2X2 inst_cellmath__43_0_I541 (.Y(N2618), .A(N3391), .B(N9379));
NOR2X4 inst_cellmath__43_0_I542 (.Y(N3544), .A(N2849), .B(N9379));
NOR2X4 inst_cellmath__43_0_I543 (.Y(N2352), .A(N2317), .B(N9379));
INVXL inst_cellmath__43_0_I544 (.Y(N3268), .A(N9379));
CLKINVX12 inst_cellmath__43_0_I545 (.Y(N3300), .A(a_man[5]));
NOR2XL inst_cellmath__43_0_I547 (.Y(N2923), .A(N3300), .B(N3614));
NOR2XL inst_cellmath__43_0_I548 (.Y(N3837), .A(N3300), .B(N3075));
NOR2XL inst_cellmath__43_0_I549 (.Y(N2653), .A(N3300), .B(N9371));
NOR2XL inst_cellmath__43_0_I550 (.Y(N3580), .A(N3300), .B(N4097));
NOR2XL inst_cellmath__43_0_I551 (.Y(N2390), .A(N3300), .B(N3571));
NOR2XL inst_cellmath__43_0_I552 (.Y(N3301), .A(N3300), .B(N3029));
NOR2XL inst_cellmath__43_0_I553 (.Y(N2120), .A(N3300), .B(N2490));
NOR2XL inst_cellmath__43_0_I554 (.Y(N3037), .A(N3300), .B(N4055));
NOR2XL inst_cellmath__43_0_I555 (.Y(N3944), .A(N3300), .B(N3526));
NOR2XL inst_cellmath__43_0_I556 (.Y(N2759), .A(N3300), .B(N2984));
NOR2XL inst_cellmath__43_0_I557 (.Y(N3687), .A(N3300), .B(N2451));
NOR2XL inst_cellmath__43_0_I558 (.Y(N2499), .A(N3300), .B(N4008));
NOR2XL inst_cellmath__43_0_I559 (.Y(N3418), .A(N3300), .B(N3479));
NOR2XL inst_cellmath__43_0_I560 (.Y(N2231), .A(N3300), .B(N2940));
NOR2XL inst_cellmath__43_0_I561 (.Y(N3146), .A(N3300), .B(N2405));
NOR2X1 inst_cellmath__43_0_I562 (.Y(N4063), .A(N3300), .B(N3963));
NOR2X1 inst_cellmath__43_0_I563 (.Y(N2880), .A(N3300), .B(N3437));
NOR2X2 inst_cellmath__43_0_I564 (.Y(N3791), .A(N3300), .B(N2895));
NOR2X1 inst_cellmath__43_0_I565 (.Y(N2609), .A(N2360), .B(N3300));
NOR2X2 inst_cellmath__43_0_I566 (.Y(N3535), .A(N3920), .B(N3300));
NOR2X1 inst_cellmath__43_0_I567 (.Y(N2344), .A(N3300), .B(N3391));
NOR2X1 inst_cellmath__43_0_I568 (.Y(N3259), .A(N3300), .B(N2849));
NOR2XL inst_cellmath__43_0_I569 (.Y(N2081), .A(N3300), .B(N2317));
INVXL inst_cellmath__43_0_I570 (.Y(N2992), .A(N3300));
CLKINVX12 inst_cellmath__43_0_I571 (.Y(N2309), .A(a_man[6]));
NOR2XL inst_cellmath__43_0_I573 (.Y(N2645), .A(N2309), .B(N3614));
NOR2XL inst_cellmath__43_0_I574 (.Y(N3567), .A(N2309), .B(N3075));
NOR2XL inst_cellmath__43_0_I575 (.Y(N2377), .A(N2309), .B(N9371));
NOR2XL inst_cellmath__43_0_I576 (.Y(N3292), .A(N2309), .B(N4097));
NOR2XL inst_cellmath__43_0_I577 (.Y(N2111), .A(N2309), .B(N3571));
NOR2XL inst_cellmath__43_0_I578 (.Y(N3025), .A(N2309), .B(N3029));
NOR2XL inst_cellmath__43_0_I579 (.Y(N3938), .A(N2309), .B(N2490));
NOR2XL inst_cellmath__43_0_I580 (.Y(N2751), .A(N2309), .B(N4055));
NOR2XL inst_cellmath__43_0_I581 (.Y(N3678), .A(N2309), .B(N3526));
NOR2XL inst_cellmath__43_0_I582 (.Y(N2488), .A(N2309), .B(N2984));
NOR2XL inst_cellmath__43_0_I583 (.Y(N3409), .A(N2309), .B(N2451));
NOR2XL inst_cellmath__43_0_I584 (.Y(N2224), .A(N2309), .B(N4008));
NOR2XL inst_cellmath__43_0_I585 (.Y(N3136), .A(N2309), .B(N3479));
NOR2XL inst_cellmath__43_0_I586 (.Y(N4051), .A(N2309), .B(N2940));
NOR2X1 inst_cellmath__43_0_I587 (.Y(N2872), .A(N2309), .B(N2405));
NOR2X1 inst_cellmath__43_0_I588 (.Y(N3781), .A(N3963), .B(N2309));
NOR2X4 inst_cellmath__43_0_I589 (.Y(N2602), .A(N2309), .B(N3437));
NOR2XL inst_cellmath__43_0_I590 (.Y(N3525), .A(N2309), .B(N2895));
NOR2X2 inst_cellmath__43_0_I591 (.Y(N2335), .A(N2309), .B(N2360));
NOR2XL inst_cellmath__43_0_I592 (.Y(N3250), .A(N2309), .B(N3920));
NOR2X1 inst_cellmath__43_0_I593 (.Y(N2073), .A(N3391), .B(N2309));
NOR2XL inst_cellmath__43_0_I594 (.Y(N2980), .A(N2309), .B(N2849));
NOR2XL inst_cellmath__43_0_I595 (.Y(N3893), .A(N2309), .B(N2317));
INVXL inst_cellmath__43_0_I596 (.Y(N2712), .A(N2309));
CLKINVX12 inst_cellmath__43_0_I597 (.Y(N3417), .A(a_man[7]));
INVX8 inst_cellmath__43_0_I4096 (.Y(N9380), .A(N3417));
INVX12 inst_cellmath__43_0_I4097 (.Y(N9381), .A(N9380));
NOR2XL inst_cellmath__43_0_I600 (.Y(N2368), .A(N9381), .B(N3614));
NOR2XL inst_cellmath__43_0_I601 (.Y(N3283), .A(N9381), .B(N3075));
NOR2XL inst_cellmath__43_0_I602 (.Y(N2102), .A(N9381), .B(N9371));
NOR2XL inst_cellmath__43_0_I603 (.Y(N3014), .A(N9381), .B(N4097));
NOR2XL inst_cellmath__43_0_I604 (.Y(N3929), .A(N9381), .B(N3571));
NOR2XL inst_cellmath__43_0_I605 (.Y(N2742), .A(N9381), .B(N3029));
NOR2XL inst_cellmath__43_0_I606 (.Y(N3671), .A(N9381), .B(N2490));
NOR2XL inst_cellmath__43_0_I607 (.Y(N2480), .A(N9381), .B(N4055));
NOR2XL inst_cellmath__43_0_I608 (.Y(N3398), .A(N9381), .B(N3526));
NOR2XL inst_cellmath__43_0_I609 (.Y(N2213), .A(N9381), .B(N2984));
NOR2XL inst_cellmath__43_0_I610 (.Y(N3128), .A(N9381), .B(N2451));
NOR2XL inst_cellmath__43_0_I611 (.Y(N4040), .A(N9381), .B(N4008));
NOR2XL inst_cellmath__43_0_I612 (.Y(N2860), .A(N9381), .B(N3479));
NOR2X1 inst_cellmath__43_0_I613 (.Y(N3774), .A(N9381), .B(N2940));
NOR2X4 inst_cellmath__43_0_I614 (.Y(N2593), .A(N2405), .B(N9381));
NOR2X2 inst_cellmath__43_0_I615 (.Y(N3514), .A(N3417), .B(N3963));
NOR2X1 inst_cellmath__43_0_I616 (.Y(N2327), .A(N3437), .B(N9381));
NOR2XL inst_cellmath__43_0_I617 (.Y(N3241), .A(N3417), .B(N2895));
NOR2XL inst_cellmath__43_0_I618 (.Y(N2066), .A(N2360), .B(N9381));
NOR2X2 inst_cellmath__43_0_I619 (.Y(N2971), .A(N3920), .B(N9381));
NOR2XL inst_cellmath__43_0_I620 (.Y(N3885), .A(N3391), .B(N9381));
NOR2XL inst_cellmath__43_0_I621 (.Y(N2705), .A(N9381), .B(N2849));
NOR2XL inst_cellmath__43_0_I622 (.Y(N3631), .A(N9381), .B(N2317));
INVXL inst_cellmath__43_0_I623 (.Y(N2438), .A(N9381));
CLKINVX12 inst_cellmath__43_0_I624 (.Y(N2878), .A(a_man[8]));
NOR2XL inst_cellmath__43_0_I626 (.Y(N2093), .A(N2878), .B(N3614));
NOR2XL inst_cellmath__43_0_I627 (.Y(N3006), .A(N2878), .B(N3075));
NOR2XL inst_cellmath__43_0_I628 (.Y(N3919), .A(N2878), .B(N9371));
NOR2XL inst_cellmath__43_0_I629 (.Y(N2734), .A(N2878), .B(N4097));
NOR2XL inst_cellmath__43_0_I630 (.Y(N3662), .A(N2878), .B(N3571));
NOR2XL inst_cellmath__43_0_I631 (.Y(N2473), .A(N2878), .B(N3029));
NOR2XL inst_cellmath__43_0_I632 (.Y(N3388), .A(N2878), .B(N2490));
NOR2XL inst_cellmath__43_0_I633 (.Y(N2205), .A(N2878), .B(N4055));
NOR2XL inst_cellmath__43_0_I634 (.Y(N3121), .A(N2878), .B(N3526));
NOR2XL inst_cellmath__43_0_I635 (.Y(N4030), .A(N2878), .B(N2984));
NOR2XL inst_cellmath__43_0_I636 (.Y(N2846), .A(N2878), .B(N2451));
NOR2XL inst_cellmath__43_0_I637 (.Y(N3764), .A(N2878), .B(N4008));
NOR2X1 inst_cellmath__43_0_I638 (.Y(N2582), .A(N3479), .B(N2878));
NOR2XL inst_cellmath__43_0_I639 (.Y(N3503), .A(N2878), .B(N2940));
NOR2X6 inst_cellmath__43_0_I640 (.Y(N2316), .A(N2878), .B(N2405));
NOR2X1 inst_cellmath__43_0_I641 (.Y(N3231), .A(N2878), .B(N3963));
NOR2X1 inst_cellmath__43_0_I642 (.Y(N2052), .A(N3437), .B(N2878));
NOR2X1 inst_cellmath__43_0_I643 (.Y(N2962), .A(N2878), .B(N2895));
NOR2X1 inst_cellmath__43_0_I644 (.Y(N3874), .A(N2360), .B(N2878));
NOR2XL inst_cellmath__43_0_I645 (.Y(N2691), .A(N2878), .B(N3920));
NOR2XL inst_cellmath__43_0_I646 (.Y(N3621), .A(N3391), .B(N2878));
NOR2XL inst_cellmath__43_0_I647 (.Y(N2430), .A(N2878), .B(N2849));
NOR2XL inst_cellmath__43_0_I648 (.Y(N3344), .A(N2878), .B(N2317));
INVXL inst_cellmath__43_0_I649 (.Y(N2167), .A(N2878));
CLKINVX8 inst_cellmath__43_0_I650 (.Y(N2342), .A(a_man[9]));
NOR2XL inst_cellmath__43_0_I652 (.Y(N3909), .A(N2342), .B(N3614));
NOR2XL inst_cellmath__43_0_I653 (.Y(N2726), .A(N2342), .B(N3075));
NOR2XL inst_cellmath__43_0_I654 (.Y(N3652), .A(N2342), .B(N9371));
NOR2XL inst_cellmath__43_0_I655 (.Y(N2465), .A(N2342), .B(N4097));
NOR2XL inst_cellmath__43_0_I656 (.Y(N3379), .A(N2342), .B(N3571));
NOR2XL inst_cellmath__43_0_I657 (.Y(N2197), .A(N2342), .B(N3029));
NOR2XL inst_cellmath__43_0_I658 (.Y(N3113), .A(N2342), .B(N2490));
NOR2XL inst_cellmath__43_0_I659 (.Y(N4021), .A(N2342), .B(N4055));
NOR2XL inst_cellmath__43_0_I660 (.Y(N2837), .A(N2342), .B(N3526));
NOR2XL inst_cellmath__43_0_I661 (.Y(N3756), .A(N2342), .B(N2984));
NOR2XL inst_cellmath__43_0_I662 (.Y(N2573), .A(N2451), .B(N2342));
NOR2X2 inst_cellmath__43_0_I663 (.Y(N3494), .A(N4008), .B(N2342));
NOR2XL inst_cellmath__43_0_I664 (.Y(N2308), .A(N3479), .B(N2342));
NOR2X2 inst_cellmath__43_0_I665 (.Y(N3224), .A(N2940), .B(N2342));
NOR2X1 inst_cellmath__43_0_I666 (.Y(N2042), .A(N2342), .B(N2405));
NOR2X2 inst_cellmath__43_0_I667 (.Y(N2955), .A(N3963), .B(N2342));
NOR2XL inst_cellmath__43_0_I668 (.Y(N3866), .A(N3437), .B(N2342));
NOR2X1 inst_cellmath__43_0_I669 (.Y(N2684), .A(N2895), .B(N2342));
NOR2XL inst_cellmath__43_0_I670 (.Y(N3612), .A(N2342), .B(N2360));
NOR2XL inst_cellmath__43_0_I671 (.Y(N2421), .A(N2342), .B(N3920));
NOR2XL inst_cellmath__43_0_I672 (.Y(N3335), .A(N2342), .B(N3391));
NOR2XL inst_cellmath__43_0_I673 (.Y(N2159), .A(N2342), .B(N2849));
NOR2XL inst_cellmath__43_0_I674 (.Y(N3070), .A(N2342), .B(N2317));
INVXL inst_cellmath__43_0_I675 (.Y(N3981), .A(N2342));
CLKINVX12 inst_cellmath__43_0_I676 (.Y(N3900), .A(a_man[10]));
NOR2XL inst_cellmath__43_0_I678 (.Y(N3642), .A(N3900), .B(N3614));
NOR2XL inst_cellmath__43_0_I679 (.Y(N2455), .A(N3900), .B(N3075));
NOR2XL inst_cellmath__43_0_I680 (.Y(N3369), .A(N3900), .B(N9371));
NOR2XL inst_cellmath__43_0_I681 (.Y(N2189), .A(N3900), .B(N4097));
NOR2XL inst_cellmath__43_0_I682 (.Y(N3104), .A(N3900), .B(N3571));
NOR2XL inst_cellmath__43_0_I683 (.Y(N4014), .A(N3900), .B(N3029));
NOR2XL inst_cellmath__43_0_I684 (.Y(N2826), .A(N3900), .B(N2490));
NOR2XL inst_cellmath__43_0_I685 (.Y(N3747), .A(N3900), .B(N4055));
NOR2XL inst_cellmath__43_0_I686 (.Y(N2563), .A(N3900), .B(N3526));
NOR2XL inst_cellmath__43_0_I687 (.Y(N3485), .A(N3900), .B(N2984));
NOR2XL inst_cellmath__43_0_I688 (.Y(N2296), .A(N3900), .B(N2451));
NOR2XL inst_cellmath__43_0_I689 (.Y(N3213), .A(N3900), .B(N4008));
NOR2X4 inst_cellmath__43_0_I690 (.Y(N2030), .A(N3479), .B(N3900));
NOR2XL inst_cellmath__43_0_I691 (.Y(N2946), .A(N3900), .B(N2940));
NOR2X4 inst_cellmath__43_0_I692 (.Y(N3854), .A(N3900), .B(N2405));
NOR2X1 inst_cellmath__43_0_I693 (.Y(N2674), .A(N3963), .B(N3900));
NOR2XL inst_cellmath__43_0_I694 (.Y(N3602), .A(N3900), .B(N3437));
NOR2XL inst_cellmath__43_0_I695 (.Y(N2411), .A(N3900), .B(N2895));
NOR2XL inst_cellmath__43_0_I696 (.Y(N3324), .A(N3900), .B(N2360));
NOR2XL inst_cellmath__43_0_I697 (.Y(N2147), .A(N3900), .B(N3920));
NOR2XL inst_cellmath__43_0_I698 (.Y(N3059), .A(N3900), .B(N3391));
NOR2XL inst_cellmath__43_0_I699 (.Y(N3969), .A(N3900), .B(N2849));
NOR2XL inst_cellmath__43_0_I700 (.Y(N2785), .A(N3900), .B(N2317));
INVXL inst_cellmath__43_0_I701 (.Y(N3710), .A(N3900));
CLKINVX8 inst_cellmath__43_0_I702 (.Y(N3370), .A(a_man[11]));
NOR2XL inst_cellmath__43_0_I704 (.Y(N3360), .A(N3370), .B(N3614));
NOR2XL inst_cellmath__43_0_I705 (.Y(N2179), .A(N3370), .B(N3075));
NOR2XL inst_cellmath__43_0_I706 (.Y(N3094), .A(N3370), .B(N9371));
NOR2XL inst_cellmath__43_0_I707 (.Y(N4005), .A(N3370), .B(N4097));
NOR2XL inst_cellmath__43_0_I708 (.Y(N2819), .A(N3370), .B(N3571));
NOR2XL inst_cellmath__43_0_I709 (.Y(N3738), .A(N3370), .B(N3029));
NOR2XL inst_cellmath__43_0_I710 (.Y(N2554), .A(N3370), .B(N2490));
NOR2XL inst_cellmath__43_0_I711 (.Y(N3472), .A(N3370), .B(N4055));
NOR2XL inst_cellmath__43_0_I712 (.Y(N2287), .A(N3370), .B(N3526));
NOR2XL inst_cellmath__43_0_I713 (.Y(N3206), .A(N3370), .B(N2984));
NOR2X2 inst_cellmath__43_0_I714 (.Y(N2022), .A(N3370), .B(N2451));
NOR2X2 inst_cellmath__43_0_I715 (.Y(N2935), .A(N4008), .B(N3370));
NOR2X1 inst_cellmath__43_0_I716 (.Y(N3847), .A(N3479), .B(N3370));
NOR2X2 inst_cellmath__43_0_I717 (.Y(N2664), .A(N2940), .B(N3370));
NOR2X2 inst_cellmath__43_0_I718 (.Y(N3594), .A(N2405), .B(N3370));
NOR2X1 inst_cellmath__43_0_I719 (.Y(N2401), .A(N3370), .B(N3963));
NOR2XL inst_cellmath__43_0_I720 (.Y(N3314), .A(N3370), .B(N3437));
NOR2XL inst_cellmath__43_0_I721 (.Y(N2135), .A(N2895), .B(N3370));
NOR2XL inst_cellmath__43_0_I722 (.Y(N3047), .A(N3370), .B(N2360));
NOR2XL inst_cellmath__43_0_I723 (.Y(N3956), .A(N3370), .B(N3920));
NOR2XL inst_cellmath__43_0_I724 (.Y(N2772), .A(N3370), .B(N3391));
NOR2XL inst_cellmath__43_0_I725 (.Y(N3698), .A(N3370), .B(N2849));
NOR2XL inst_cellmath__43_0_I726 (.Y(N2509), .A(N3370), .B(N2317));
INVXL inst_cellmath__43_0_I727 (.Y(N3432), .A(N3370));
CLKINVX8 inst_cellmath__43_0_I728 (.Y(N2828), .A(a_man[12]));
NOR2XL inst_cellmath__43_0_I730 (.Y(N3085), .A(N2828), .B(N3614));
NOR2XL inst_cellmath__43_0_I731 (.Y(N3998), .A(N2828), .B(N3075));
NOR2XL inst_cellmath__43_0_I732 (.Y(N2810), .A(N2828), .B(N9371));
NOR2XL inst_cellmath__43_0_I733 (.Y(N3730), .A(N2828), .B(N4097));
NOR2XL inst_cellmath__43_0_I734 (.Y(N2547), .A(N2828), .B(N3571));
NOR2XL inst_cellmath__43_0_I735 (.Y(N3463), .A(N2828), .B(N3029));
NOR2XL inst_cellmath__43_0_I736 (.Y(N2278), .A(N2828), .B(N2490));
NOR2XL inst_cellmath__43_0_I737 (.Y(N3198), .A(N2828), .B(N4055));
NOR2XL inst_cellmath__43_0_I738 (.Y(N2013), .A(N2828), .B(N3526));
NOR2X2 inst_cellmath__43_0_I739 (.Y(N2926), .A(N2984), .B(N2828));
NOR2X4 inst_cellmath__43_0_I740 (.Y(N3839), .A(N2451), .B(N2828));
NOR2X1 inst_cellmath__43_0_I741 (.Y(N2655), .A(N4008), .B(N2828));
NOR2X2 inst_cellmath__43_0_I742 (.Y(N3583), .A(N2828), .B(N3479));
NOR2XL inst_cellmath__43_0_I743 (.Y(N2393), .A(N2940), .B(N2828));
NOR2X1 inst_cellmath__43_0_I744 (.Y(N3304), .A(N2828), .B(N2405));
NOR2XL inst_cellmath__43_0_I745 (.Y(N2123), .A(N2828), .B(N3963));
NOR2XL inst_cellmath__43_0_I746 (.Y(N3040), .A(N2828), .B(N3437));
NOR2XL inst_cellmath__43_0_I747 (.Y(N3947), .A(N2828), .B(N2895));
NOR2XL inst_cellmath__43_0_I748 (.Y(N2762), .A(N2828), .B(N2360));
NOR2XL inst_cellmath__43_0_I749 (.Y(N3690), .A(N2828), .B(N3920));
NOR2XL inst_cellmath__43_0_I750 (.Y(N2503), .A(N2828), .B(N3391));
NOR2XL inst_cellmath__43_0_I751 (.Y(N3423), .A(N2828), .B(N2849));
NOR2XL inst_cellmath__43_0_I752 (.Y(N2234), .A(N2828), .B(N2317));
INVXL inst_cellmath__43_0_I753 (.Y(N3150), .A(N2828));
CLKINVX12 inst_cellmath__43_0_I754 (.Y(N2297), .A(a_man[13]));
NOR2XL inst_cellmath__43_0_I756 (.Y(N2800), .A(N2297), .B(N3614));
NOR2XL inst_cellmath__43_0_I757 (.Y(N3721), .A(N2297), .B(N3075));
NOR2XL inst_cellmath__43_0_I758 (.Y(N2537), .A(N2297), .B(N9371));
NOR2XL inst_cellmath__43_0_I759 (.Y(N3456), .A(N2297), .B(N4097));
NOR2XL inst_cellmath__43_0_I760 (.Y(N2265), .A(N2297), .B(N3571));
NOR2XL inst_cellmath__43_0_I761 (.Y(N3190), .A(N2297), .B(N3029));
NOR2XL inst_cellmath__43_0_I762 (.Y(N4100), .A(N2297), .B(N2490));
NOR2XL inst_cellmath__43_0_I763 (.Y(N2914), .A(N2297), .B(N4055));
NOR2X1 inst_cellmath__43_0_I764 (.Y(N3830), .A(N3526), .B(N2297));
NOR2X1 inst_cellmath__43_0_I765 (.Y(N2648), .A(N2984), .B(N2297));
NOR2X1 inst_cellmath__43_0_I766 (.Y(N3572), .A(N2297), .B(N2451));
NOR2X1 inst_cellmath__43_0_I767 (.Y(N2383), .A(N2297), .B(N4008));
NOR2X1 inst_cellmath__43_0_I768 (.Y(N3295), .A(N2297), .B(N3479));
NOR2XL inst_cellmath__43_0_I769 (.Y(N2115), .A(N2297), .B(N2940));
NOR2XL inst_cellmath__43_0_I770 (.Y(N3032), .A(N2297), .B(N2405));
NOR2XL inst_cellmath__43_0_I771 (.Y(N3941), .A(N2297), .B(N3963));
NOR2XL inst_cellmath__43_0_I772 (.Y(N2755), .A(N2297), .B(N3437));
NOR2XL inst_cellmath__43_0_I773 (.Y(N3684), .A(N2297), .B(N2895));
NOR2XL inst_cellmath__43_0_I774 (.Y(N2493), .A(N2297), .B(N2360));
NOR2XL inst_cellmath__43_0_I775 (.Y(N3413), .A(N2297), .B(N3920));
NOR2XL inst_cellmath__43_0_I776 (.Y(N2227), .A(N2297), .B(N3391));
NOR2XL inst_cellmath__43_0_I777 (.Y(N3142), .A(N2297), .B(N2849));
NOR2XL inst_cellmath__43_0_I778 (.Y(N4056), .A(N2297), .B(N2317));
INVXL inst_cellmath__43_0_I779 (.Y(N2876), .A(N2297));
CLKINVX6 inst_cellmath__43_0_I780 (.Y(N3856), .A(a_man[14]));
NOR2XL inst_cellmath__43_0_I782 (.Y(N2528), .A(N3856), .B(N3614));
NOR2XL inst_cellmath__43_0_I783 (.Y(N3448), .A(N3856), .B(N3075));
NOR2XL inst_cellmath__43_0_I784 (.Y(N2255), .A(N3856), .B(N9371));
NOR2XL inst_cellmath__43_0_I785 (.Y(N3179), .A(N3856), .B(N4097));
NOR2XL inst_cellmath__43_0_I786 (.Y(N4089), .A(N3856), .B(N3571));
NOR2XL inst_cellmath__43_0_I787 (.Y(N2905), .A(N3029), .B(N3856));
NOR2XL inst_cellmath__43_0_I788 (.Y(N3820), .A(N3856), .B(N2490));
NOR2XL inst_cellmath__43_0_I789 (.Y(N2638), .A(N3856), .B(N4055));
NOR2X4 inst_cellmath__43_0_I790 (.Y(N3561), .A(N3526), .B(N3856));
NOR2X1 inst_cellmath__43_0_I791 (.Y(N2373), .A(N2984), .B(N3856));
NOR2X1 inst_cellmath__43_0_I792 (.Y(N3286), .A(N3856), .B(N2451));
NOR2X2 inst_cellmath__43_0_I793 (.Y(N2105), .A(N4008), .B(N3856));
NOR2X1 inst_cellmath__43_0_I794 (.Y(N3020), .A(N3856), .B(N3479));
NOR2XL inst_cellmath__43_0_I795 (.Y(N3932), .A(N3856), .B(N2940));
NOR2XL inst_cellmath__43_0_I796 (.Y(N2746), .A(N3856), .B(N2405));
NOR2XL inst_cellmath__43_0_I797 (.Y(N3676), .A(N3856), .B(N3963));
NOR2XL inst_cellmath__43_0_I798 (.Y(N2484), .A(N3856), .B(N3437));
NOR2XL inst_cellmath__43_0_I799 (.Y(N3401), .A(N3856), .B(N2895));
NOR2XL inst_cellmath__43_0_I800 (.Y(N2218), .A(N3856), .B(N2360));
NOR2XL inst_cellmath__43_0_I801 (.Y(N3131), .A(N3856), .B(N3920));
NOR2XL inst_cellmath__43_0_I802 (.Y(N4045), .A(N3856), .B(N3391));
NOR2XL inst_cellmath__43_0_I803 (.Y(N2867), .A(N3856), .B(N2849));
NOR2XL inst_cellmath__43_0_I804 (.Y(N3777), .A(N3856), .B(N2317));
INVXL inst_cellmath__43_0_I805 (.Y(N2597), .A(N3856));
CLKINVX8 inst_cellmath__43_0_I806 (.Y(N3328), .A(a_man[15]));
NOR2XL inst_cellmath__43_0_I808 (.Y(N2246), .A(N3328), .B(N3614));
NOR2XL inst_cellmath__43_0_I809 (.Y(N3166), .A(N3328), .B(N3075));
NOR2XL inst_cellmath__43_0_I810 (.Y(N4082), .A(N3328), .B(N9371));
NOR2XL inst_cellmath__43_0_I811 (.Y(N2897), .A(N3328), .B(N4097));
NOR2XL inst_cellmath__43_0_I812 (.Y(N3808), .A(N3328), .B(N3571));
NOR2XL inst_cellmath__43_0_I813 (.Y(N2630), .A(N3029), .B(N3328));
NOR2XL inst_cellmath__43_0_I814 (.Y(N3552), .A(N2490), .B(N3328));
NOR2X4 inst_cellmath__43_0_I815 (.Y(N2363), .A(N4055), .B(N3328));
NOR2XL inst_cellmath__43_0_I816 (.Y(N3279), .A(N3328), .B(N3526));
NOR2X2 inst_cellmath__43_0_I817 (.Y(N2095), .A(N3328), .B(N2984));
NOR2XL inst_cellmath__43_0_I818 (.Y(N3010), .A(N3328), .B(N2451));
NOR2X1 inst_cellmath__43_0_I819 (.Y(N3922), .A(N3328), .B(N4008));
NOR2XL inst_cellmath__43_0_I820 (.Y(N2736), .A(N3328), .B(N3479));
NOR2XL inst_cellmath__43_0_I821 (.Y(N3668), .A(N3328), .B(N2940));
NOR2X1 inst_cellmath__43_0_I822 (.Y(N2475), .A(N2405), .B(N3328));
NOR2XL inst_cellmath__43_0_I823 (.Y(N3392), .A(N3328), .B(N3963));
NOR2XL inst_cellmath__43_0_I824 (.Y(N2210), .A(N3328), .B(N3437));
NOR2XL inst_cellmath__43_0_I825 (.Y(N3123), .A(N3328), .B(N2895));
NOR2XL inst_cellmath__43_0_I826 (.Y(N4033), .A(N3328), .B(N2360));
NOR2XL inst_cellmath__43_0_I827 (.Y(N2853), .A(N3328), .B(N3920));
NOR2XL inst_cellmath__43_0_I828 (.Y(N3766), .A(N3328), .B(N3391));
NOR2XL inst_cellmath__43_0_I829 (.Y(N2585), .A(N3328), .B(N2849));
NOR2XL inst_cellmath__43_0_I830 (.Y(N3508), .A(N3328), .B(N2317));
INVXL inst_cellmath__43_0_I831 (.Y(N2319), .A(N3328));
CLKINVX12 inst_cellmath__43_0_I832 (.Y(N2786), .A(a_man[16]));
NOR2XL inst_cellmath__43_0_I833 (.Y(N4072), .A(N2786), .B(N3614));
NOR2XL inst_cellmath__43_0_I834 (.Y(N2887), .A(N2786), .B(N3075));
NOR2XL inst_cellmath__43_0_I835 (.Y(N3799), .A(N2786), .B(N9371));
NOR2XL inst_cellmath__43_0_I836 (.Y(N2621), .A(N2786), .B(N4097));
NOR2XL inst_cellmath__43_0_I837 (.Y(N3543), .A(N2786), .B(N3571));
NOR2XL inst_cellmath__43_0_I838 (.Y(N2351), .A(N2786), .B(N3029));
NOR2X2 inst_cellmath__43_0_I839 (.Y(N3271), .A(N2786), .B(N2490));
NOR2X1 inst_cellmath__43_0_I840 (.Y(N2088), .A(N2786), .B(N4055));
NOR2X2 inst_cellmath__43_0_I841 (.Y(N3000), .A(N3526), .B(N2786));
NOR2X2 inst_cellmath__43_0_I842 (.Y(N3913), .A(N2984), .B(N2786));
NOR2XL inst_cellmath__43_0_I843 (.Y(N2729), .A(N2786), .B(N2451));
NOR2XL inst_cellmath__43_0_I844 (.Y(N3655), .A(N2786), .B(N4008));
NOR2XL inst_cellmath__43_0_I845 (.Y(N2469), .A(N2786), .B(N3479));
NOR2XL inst_cellmath__43_0_I846 (.Y(N3383), .A(N2786), .B(N2940));
NOR2X1 inst_cellmath__43_0_I847 (.Y(N2200), .A(N2786), .B(N2405));
NOR2XL inst_cellmath__43_0_I848 (.Y(N3117), .A(N2786), .B(N3963));
NOR2XL inst_cellmath__43_0_I849 (.Y(N4024), .A(N2786), .B(N3437));
NOR2XL inst_cellmath__43_0_I850 (.Y(N2842), .A(N2786), .B(N2895));
NOR2XL inst_cellmath__43_0_I851 (.Y(N3758), .A(N2786), .B(N2360));
NOR2XL inst_cellmath__43_0_I852 (.Y(N2575), .A(N2786), .B(N3920));
NOR2XL inst_cellmath__43_0_I853 (.Y(N3499), .A(N2786), .B(N3391));
NOR2XL inst_cellmath__43_0_I854 (.Y(N2311), .A(N2786), .B(N2849));
NOR2XL inst_cellmath__43_0_I855 (.Y(N3226), .A(N2786), .B(N2317));
INVXL inst_cellmath__43_0_I856 (.Y(N2047), .A(N2786));
CLKINVX6 inst_cellmath__43_0_I857 (.Y(N2251), .A(a_man[17]));
NOR2XL inst_cellmath__43_0_I858 (.Y(N3790), .A(N2251), .B(N3614));
NOR2XL inst_cellmath__43_0_I859 (.Y(N2612), .A(N2251), .B(N3075));
NOR2XL inst_cellmath__43_0_I860 (.Y(N3534), .A(N2251), .B(N9371));
NOR2XL inst_cellmath__43_0_I861 (.Y(N2343), .A(N2251), .B(N4097));
NOR2XL inst_cellmath__43_0_I862 (.Y(N3262), .A(N3571), .B(N2251));
NOR2X1 inst_cellmath__43_0_I863 (.Y(N2080), .A(N3029), .B(N2251));
NOR2X1 inst_cellmath__43_0_I864 (.Y(N2991), .A(N2490), .B(N2251));
NOR2X1 inst_cellmath__43_0_I865 (.Y(N3904), .A(N4055), .B(N2251));
NOR2X2 inst_cellmath__43_0_I866 (.Y(N2720), .A(N2251), .B(N3526));
NOR2XL inst_cellmath__43_0_I867 (.Y(N3644), .A(N2251), .B(N2984));
NOR2XL inst_cellmath__43_0_I868 (.Y(N2461), .A(N2251), .B(N2451));
NOR2XL inst_cellmath__43_0_I869 (.Y(N3373), .A(N2251), .B(N4008));
NOR2XL inst_cellmath__43_0_I870 (.Y(N2191), .A(N2251), .B(N3479));
NOR2XL inst_cellmath__43_0_I871 (.Y(N3108), .A(N2251), .B(N2940));
NOR2XL inst_cellmath__43_0_I872 (.Y(N4017), .A(N2251), .B(N2405));
NOR2XL inst_cellmath__43_0_I873 (.Y(N2829), .A(N2251), .B(N3963));
NOR2XL inst_cellmath__43_0_I874 (.Y(N3751), .A(N2251), .B(N3437));
NOR2XL inst_cellmath__43_0_I875 (.Y(N2567), .A(N2251), .B(N2895));
NOR2XL inst_cellmath__43_0_I876 (.Y(N3487), .A(N2251), .B(N2360));
NOR2XL inst_cellmath__43_0_I877 (.Y(N2301), .A(N2251), .B(N3920));
NOR2XL inst_cellmath__43_0_I878 (.Y(N3216), .A(N2251), .B(N3391));
NOR2XL inst_cellmath__43_0_I879 (.Y(N2034), .A(N2251), .B(N2849));
NOR2XL inst_cellmath__43_0_I880 (.Y(N2950), .A(N2251), .B(N2317));
INVXL inst_cellmath__43_0_I881 (.Y(N3858), .A(N2251));
CLKINVX6 inst_cellmath__43_0_I882 (.Y(N3361), .A(a_man[18]));
NOR2XL inst_cellmath__43_0_I883 (.Y(N3524), .A(N3361), .B(N3614));
NOR2XL inst_cellmath__43_0_I884 (.Y(N2334), .A(N3361), .B(N3075));
NOR2X1 inst_cellmath__43_0_I885 (.Y(N3253), .A(N3361), .B(N9371));
NOR2X1 inst_cellmath__43_0_I886 (.Y(N2072), .A(N4097), .B(N3361));
NOR2X1 inst_cellmath__43_0_I887 (.Y(N2979), .A(N3571), .B(N3361));
NOR2XL inst_cellmath__43_0_I888 (.Y(N3896), .A(N3361), .B(N3029));
NOR2X2 inst_cellmath__43_0_I889 (.Y(N2711), .A(N3361), .B(N2490));
NOR2X1 inst_cellmath__43_0_I890 (.Y(N3637), .A(N3361), .B(N4055));
NOR2XL inst_cellmath__43_0_I891 (.Y(N2450), .A(N3361), .B(N3526));
NOR2XL inst_cellmath__43_0_I892 (.Y(N3364), .A(N3361), .B(N2984));
NOR2XL inst_cellmath__43_0_I893 (.Y(N2182), .A(N3361), .B(N2451));
NOR2XL inst_cellmath__43_0_I894 (.Y(N3099), .A(N3361), .B(N4008));
NOR2XL inst_cellmath__43_0_I895 (.Y(N4007), .A(N3361), .B(N3479));
NOR2XL inst_cellmath__43_0_I896 (.Y(N2821), .A(N3361), .B(N2940));
NOR2X1 inst_cellmath__43_0_I897 (.Y(N3743), .A(N2405), .B(N3361));
NOR2XL inst_cellmath__43_0_I898 (.Y(N2556), .A(N3361), .B(N3963));
NOR2XL inst_cellmath__43_0_I899 (.Y(N3475), .A(N3361), .B(N3437));
NOR2XL inst_cellmath__43_0_I900 (.Y(N2291), .A(N3361), .B(N2895));
NOR2XL inst_cellmath__43_0_I901 (.Y(N3208), .A(N3361), .B(N2360));
NOR2XL inst_cellmath__43_0_I902 (.Y(N2024), .A(N3361), .B(N3920));
NOR2XL inst_cellmath__43_0_I903 (.Y(N2939), .A(N3361), .B(N3391));
NOR2XL inst_cellmath__43_0_I904 (.Y(N3849), .A(N3361), .B(N2849));
NOR2XL inst_cellmath__43_0_I905 (.Y(N2667), .A(N3361), .B(N2317));
INVXL inst_cellmath__43_0_I906 (.Y(N3597), .A(N3361));
CLKINVX4 inst_cellmath__43_0_I907 (.Y(N2367), .A(a_man[19]));
NOR2XL inst_cellmath__43_0_I908 (.Y(N3240), .A(N2367), .B(N3614));
NOR2XL inst_cellmath__43_0_I909 (.Y(N2065), .A(N2367), .B(N3075));
NOR2XL inst_cellmath__43_0_I910 (.Y(N2970), .A(N2367), .B(N1902));
NOR2XL inst_cellmath__43_0_I911 (.Y(N3888), .A(N2367), .B(N4097));
NOR2XL inst_cellmath__43_0_I912 (.Y(N2704), .A(N2367), .B(N3571));
NOR2XL inst_cellmath__43_0_I913 (.Y(N3630), .A(N2367), .B(N3029));
NOR2XL inst_cellmath__43_0_I914 (.Y(N2441), .A(N2367), .B(N2490));
NOR2XL inst_cellmath__43_0_I915 (.Y(N3355), .A(N2367), .B(N4055));
NOR2XL inst_cellmath__43_0_I916 (.Y(N2174), .A(N2367), .B(N3526));
NOR2XL inst_cellmath__43_0_I917 (.Y(N3091), .A(N2367), .B(N2984));
NOR2XL inst_cellmath__43_0_I918 (.Y(N4001), .A(N2367), .B(N2451));
NOR2XL inst_cellmath__43_0_I919 (.Y(N2814), .A(N2367), .B(N4008));
NOR2XL inst_cellmath__43_0_I920 (.Y(N3735), .A(N2367), .B(N3479));
NOR2XL inst_cellmath__43_0_I921 (.Y(N2550), .A(N2367), .B(N2940));
NOR2XL inst_cellmath__43_0_I922 (.Y(N3468), .A(N2367), .B(N2405));
NOR2XL inst_cellmath__43_0_I923 (.Y(N2284), .A(N2367), .B(N3963));
NOR2XL inst_cellmath__43_0_I924 (.Y(N3201), .A(N2367), .B(N3437));
NOR2XL inst_cellmath__43_0_I925 (.Y(N2016), .A(N2367), .B(N2895));
NOR2XL inst_cellmath__43_0_I926 (.Y(N2930), .A(N2367), .B(N2360));
NOR2XL inst_cellmath__43_0_I927 (.Y(N3842), .A(N2367), .B(N3920));
NOR2XL inst_cellmath__43_0_I928 (.Y(N2658), .A(N2367), .B(N3391));
NOR2XL inst_cellmath__43_0_I929 (.Y(N3587), .A(N2367), .B(N2849));
NOR2XL inst_cellmath__43_0_I930 (.Y(N2396), .A(N2367), .B(N2317));
INVXL inst_cellmath__43_0_I931 (.Y(N3308), .A(N2367));
CLKINVX8 inst_cellmath__43_0_I932 (.Y(N3927), .A(a_man[20]));
NOR2XL inst_cellmath__43_0_I934 (.Y(N2961), .A(N3927), .B(N3614));
NOR2XL inst_cellmath__43_0_I935 (.Y(N3873), .A(N3927), .B(N3075));
NOR2XL inst_cellmath__43_0_I936 (.Y(N2693), .A(N3927), .B(N9371));
NOR2XL inst_cellmath__43_0_I937 (.Y(N3620), .A(N3927), .B(N4097));
NOR2X2 inst_cellmath__43_0_I938 (.Y(N2429), .A(N3927), .B(N3571));
NOR2XL inst_cellmath__43_0_I939 (.Y(N3346), .A(N3927), .B(N3029));
NOR2XL inst_cellmath__43_0_I940 (.Y(N2166), .A(N3927), .B(N2490));
NOR2XL inst_cellmath__43_0_I941 (.Y(N3080), .A(N3927), .B(N4055));
NOR2XL inst_cellmath__43_0_I942 (.Y(N3991), .A(N3927), .B(N3526));
NOR2XL inst_cellmath__43_0_I943 (.Y(N2805), .A(N3927), .B(N2984));
NOR2XL inst_cellmath__43_0_I944 (.Y(N3727), .A(N3927), .B(N2451));
NOR2XL inst_cellmath__43_0_I945 (.Y(N2540), .A(N3927), .B(N4008));
NOR2XL inst_cellmath__43_0_I946 (.Y(N3459), .A(N3927), .B(N3479));
NOR2XL inst_cellmath__43_0_I947 (.Y(N2273), .A(N3927), .B(N2940));
NOR2XL inst_cellmath__43_0_I948 (.Y(N3192), .A(N3927), .B(N2405));
NOR2XL inst_cellmath__43_0_I949 (.Y(N4104), .A(N3927), .B(N3963));
NOR2XL inst_cellmath__43_0_I950 (.Y(N2920), .A(N3927), .B(N3437));
NOR2XL inst_cellmath__43_0_I951 (.Y(N3832), .A(N3927), .B(N2895));
NOR2XL inst_cellmath__43_0_I952 (.Y(N2650), .A(N3927), .B(N2360));
NOR2XL inst_cellmath__43_0_I953 (.Y(N3578), .A(N3927), .B(N3920));
NOR2XL inst_cellmath__43_0_I954 (.Y(N2386), .A(N3927), .B(N3391));
NOR2XL inst_cellmath__43_0_I955 (.Y(N3298), .A(N3927), .B(N2849));
NOR2XL inst_cellmath__43_0_I956 (.Y(N2119), .A(N3927), .B(N2317));
INVXL inst_cellmath__43_0_I957 (.Y(N3035), .A(N3927));
CLKINVX6 inst_cellmath__43_0_I958 (.Y(N3397), .A(a_man[21]));
NOR2XL inst_cellmath__43_0_I959 (.Y(N2686), .A(N3397), .B(N3614));
NOR2XL inst_cellmath__43_0_I960 (.Y(N3611), .A(N3397), .B(N3075));
NOR2XL inst_cellmath__43_0_I961 (.Y(N2420), .A(N3397), .B(N9371));
NOR2X1 inst_cellmath__43_0_I962 (.Y(N3337), .A(N3397), .B(N4097));
NOR2XL inst_cellmath__43_0_I963 (.Y(N2158), .A(N3397), .B(N3571));
NOR2XL inst_cellmath__43_0_I964 (.Y(N3069), .A(N3397), .B(N3029));
NOR2XL inst_cellmath__43_0_I965 (.Y(N3983), .A(N3397), .B(N2490));
NOR2XL inst_cellmath__43_0_I966 (.Y(N2795), .A(N3397), .B(N4055));
NOR2XL inst_cellmath__43_0_I967 (.Y(N3717), .A(N3397), .B(N3526));
NOR2XL inst_cellmath__43_0_I968 (.Y(N2530), .A(N3397), .B(N2984));
NOR2XL inst_cellmath__43_0_I969 (.Y(N3452), .A(N3397), .B(N2451));
NOR2XL inst_cellmath__43_0_I970 (.Y(N2259), .A(N3397), .B(N4008));
NOR2XL inst_cellmath__43_0_I971 (.Y(N3183), .A(N3397), .B(N3479));
NOR2XL inst_cellmath__43_0_I972 (.Y(N4094), .A(N3397), .B(N2940));
NOR2XL inst_cellmath__43_0_I973 (.Y(N2909), .A(N3397), .B(N2405));
NOR2XL inst_cellmath__43_0_I974 (.Y(N3824), .A(N3397), .B(N3963));
NOR2XL inst_cellmath__43_0_I975 (.Y(N2642), .A(N3397), .B(N3437));
NOR2XL inst_cellmath__43_0_I976 (.Y(N3565), .A(N3397), .B(N2895));
NOR2XL inst_cellmath__43_0_I977 (.Y(N2375), .A(N3397), .B(N2360));
NOR2XL inst_cellmath__43_0_I978 (.Y(N3288), .A(N3397), .B(N3920));
NOR2XL inst_cellmath__43_0_I979 (.Y(N2110), .A(N3397), .B(N3391));
NOR2XL inst_cellmath__43_0_I980 (.Y(N3023), .A(N3397), .B(N2849));
NOR2XL inst_cellmath__43_0_I981 (.Y(N3934), .A(N3397), .B(N2317));
INVXL inst_cellmath__43_0_I982 (.Y(N2750), .A(N3397));
CLKINVX8 inst_cellmath__43_0_I983 (.Y(N2857), .A(a_man[22]));
NOR2XL inst_cellmath__43_0_I984 (.Y(N2410), .A(N2857), .B(N3614));
NOR2XL inst_cellmath__43_0_I985 (.Y(N3327), .A(N2857), .B(N3075));
NOR2X2 inst_cellmath__43_0_I986 (.Y(N2146), .A(N2857), .B(N1902));
NOR2XL inst_cellmath__43_0_I987 (.Y(N3058), .A(N2857), .B(N4097));
NOR2XL inst_cellmath__43_0_I988 (.Y(N3972), .A(N2857), .B(N3571));
NOR2XL inst_cellmath__43_0_I989 (.Y(N2784), .A(N2857), .B(N3029));
NOR2XL inst_cellmath__43_0_I990 (.Y(N3709), .A(N2857), .B(N2490));
NOR2XL inst_cellmath__43_0_I991 (.Y(N2521), .A(N2857), .B(N4055));
NOR2XL inst_cellmath__43_0_I992 (.Y(N3444), .A(N2857), .B(N3526));
NOR2XL inst_cellmath__43_0_I993 (.Y(N2249), .A(N2857), .B(N2984));
NOR2XL inst_cellmath__43_0_I994 (.Y(N3172), .A(N2857), .B(N2451));
NOR2XL inst_cellmath__43_0_I995 (.Y(N4084), .A(N2857), .B(N4008));
NOR2XL inst_cellmath__43_0_I996 (.Y(N2901), .A(N2857), .B(N3479));
NOR2XL inst_cellmath__43_0_I997 (.Y(N3814), .A(N2857), .B(N2940));
NOR2XL inst_cellmath__43_0_I998 (.Y(N2633), .A(N2857), .B(N2405));
NOR2XL inst_cellmath__43_0_I999 (.Y(N3556), .A(N2857), .B(N3963));
NOR2XL inst_cellmath__43_0_I1000 (.Y(N2366), .A(N2857), .B(N3437));
NOR2XL inst_cellmath__43_0_I1001 (.Y(N3281), .A(N2857), .B(N2895));
NOR2XL inst_cellmath__43_0_I1002 (.Y(N2099), .A(N2857), .B(N2360));
NOR2XL inst_cellmath__43_0_I1003 (.Y(N3012), .A(N2857), .B(N3920));
NOR2XL inst_cellmath__43_0_I1004 (.Y(N3926), .A(N2857), .B(N3391));
NOR2XL inst_cellmath__43_0_I1005 (.Y(N2740), .A(N2857), .B(N2849));
NOR2XL inst_cellmath__43_0_I1006 (.Y(N3670), .A(N2857), .B(N2317));
INVXL inst_cellmath__43_0_I1007 (.Y(N2478), .A(N2857));
INVX1 inst_cellmath__43_0_I1008 (.Y(N2400), .A(N3614));
INVXL inst_cellmath__43_0_I1009 (.Y(N3317), .A(N3075));
CLKINVX4 inst_cellmath__43_0_I1010 (.Y(N2134), .A(N9371));
INVXL inst_cellmath__43_0_I1011 (.Y(N3046), .A(N4097));
INVXL inst_cellmath__43_0_I1012 (.Y(N3959), .A(N3571));
INVXL inst_cellmath__43_0_I1013 (.Y(N2771), .A(N3029));
INVXL inst_cellmath__43_0_I1014 (.Y(N3697), .A(N2490));
INVXL inst_cellmath__43_0_I1015 (.Y(N2512), .A(N4055));
INVXL inst_cellmath__43_0_I1016 (.Y(N3431), .A(N3526));
INVXL inst_cellmath__43_0_I1017 (.Y(N2239), .A(N2984));
INVXL inst_cellmath__43_0_I1018 (.Y(N3162), .A(N2451));
INVXL inst_cellmath__43_0_I1019 (.Y(N4075), .A(N4008));
INVXL inst_cellmath__43_0_I1020 (.Y(N2890), .A(N3479));
INVXL inst_cellmath__43_0_I1021 (.Y(N3805), .A(N2940));
INVXL inst_cellmath__43_0_I1022 (.Y(N2623), .A(N2405));
INVXL inst_cellmath__43_0_I1023 (.Y(N3546), .A(N3963));
INVXL inst_cellmath__43_0_I1024 (.Y(N2357), .A(N3437));
INVXL inst_cellmath__43_0_I1025 (.Y(N3274), .A(N2895));
INVXL inst_cellmath__43_0_I1026 (.Y(N2090), .A(N2360));
INVXL inst_cellmath__43_0_I1027 (.Y(N3005), .A(N3920));
INVXL inst_cellmath__43_0_I1028 (.Y(N3915), .A(N3391));
INVXL inst_cellmath__43_0_I1029 (.Y(N2731), .A(N2849));
INVXL inst_cellmath__43_0_I1030 (.Y(N3661), .A(N2317));
ADDHX1 inst_cellmath__43_0_I1031 (.CO(N2882), .S(N2428), .A(N4036), .B(N2843));
ADDHX1 inst_cellmath__43_0_I1032 (.CO(N3796), .S(N3342), .A(N2855), .B(N3760));
ADDFX1 inst_cellmath__43_0_I1033 (.CO(N2614), .S(N2162), .A(N3480), .B(N2570), .CI(N2882));
ADDHX1 inst_cellmath__43_0_I1034 (.CO(N3537), .S(N3079), .A(N3769), .B(N2578));
ADDFXL inst_cellmath__43_0_I1035 (.CO(N2348), .S(N3988), .A(N2292), .B(N3491), .CI(N3203));
ADDFX1 inst_cellmath__43_0_I1036 (.CO(N3264), .S(N2799), .A(N3079), .B(N3796), .CI(N3988));
ADDHX1 inst_cellmath__43_0_I1037 (.CO(N2083), .S(N3724), .A(N2589), .B(N3501));
ADDFX1 inst_cellmath__43_0_I1038 (.CO(N2996), .S(N2536), .A(N3211), .B(N2302), .CI(N2019));
ADDFX1 inst_cellmath__43_0_I1039 (.CO(N3906), .S(N3455), .A(N3537), .B(N2923), .CI(N3724));
ADDFX1 inst_cellmath__43_0_I1040 (.CO(N2722), .S(N2269), .A(N2536), .B(N2348), .CI(N3264));
ADDHX1 inst_cellmath__43_0_I1041 (.CO(N3650), .S(N3189), .A(N3511), .B(N2313));
ADDFX1 inst_cellmath__43_0_I1042 (.CO(N2463), .S(N4099), .A(N2027), .B(N3220), .CI(N2932));
ADDFX1 inst_cellmath__43_0_I1043 (.CO(N3375), .S(N2916), .A(N2645), .B(N3837), .CI(N2083));
ADDFX1 inst_cellmath__43_0_I1044 (.CO(N2196), .S(N3829), .A(N2996), .B(N3189), .CI(N4099));
ADDFX1 inst_cellmath__43_0_I1045 (.CO(N3110), .S(N2647), .A(N2916), .B(N3906), .CI(N3829));
ADDHX1 inst_cellmath__43_0_I1046 (.CO(N4019), .S(N3575), .A(N2323), .B(N3229));
ADDFX1 inst_cellmath__43_0_I1047 (.CO(N2835), .S(N2382), .A(N2941), .B(N2038), .CI(N3844));
ADDFX1 inst_cellmath__43_0_I1048 (.CO(N3754), .S(N3294), .A(N3567), .B(N2653), .CI(N2368));
ADDFX1 inst_cellmath__43_0_I1049 (.CO(N2569), .S(N2117), .A(N3575), .B(N3650), .CI(N2463));
ADDFX1 inst_cellmath__43_0_I1050 (.CO(N3493), .S(N3031), .A(N3294), .B(N2382), .CI(N3375));
ADDFX1 inst_cellmath__43_0_I1051 (.CO(N2304), .S(N3940), .A(N2117), .B(N2196), .CI(N3031));
ADDHX1 inst_cellmath__43_0_I1052 (.CO(N3219), .S(N2757), .A(N3236), .B(N2048));
ADDFX1 inst_cellmath__43_0_I1053 (.CO(N2041), .S(N3683), .A(N3852), .B(N2951), .CI(N2661));
ADDFX1 inst_cellmath__43_0_I1054 (.CO(N2953), .S(N2492), .A(N3580), .B(N2377), .CI(N3283));
ADDFX1 inst_cellmath__43_0_I1055 (.CO(N3862), .S(N3415), .A(N4019), .B(N2093), .CI(N2757));
ADDFX1 inst_cellmath__43_0_I1056 (.CO(N2682), .S(N2226), .A(N3754), .B(N2835), .CI(N3683));
ADDFX1 inst_cellmath__43_0_I1057 (.CO(N3608), .S(N3141), .A(N2569), .B(N2492), .CI(N3415));
ADDFX1 inst_cellmath__43_0_I1058 (.CO(N2417), .S(N4059), .A(N2226), .B(N3493), .CI(N3141));
ADDHX1 inst_cellmath__43_0_I1059 (.CO(N3334), .S(N2875), .A(N2059), .B(N2959));
ADDFX1 inst_cellmath__43_0_I1060 (.CO(N2154), .S(N3786), .A(N2671), .B(N3863), .CI(N3589));
ADDFX1 inst_cellmath__43_0_I1061 (.CO(N3065), .S(N2607), .A(N3292), .B(N2390), .CI(N2102));
ADDFX1 inst_cellmath__43_0_I1062 (.CO(N3978), .S(N3529), .A(N3909), .B(N3006), .CI(N3219));
ADDFXL inst_cellmath__43_0_I1063 (.CO(N2790), .S(N2339), .A(N2875), .B(N2041), .CI(N2953));
ADDFX1 inst_cellmath__43_0_I1064 (.CO(N3714), .S(N3256), .A(N2607), .B(N3786), .CI(N3862));
ADDFXL inst_cellmath__43_0_I1065 (.CO(N2527), .S(N2077), .A(N2682), .B(N3529), .CI(N2339));
ADDFX1 inst_cellmath__43_0_I1066 (.CO(N3447), .S(N2987), .A(N3256), .B(N3608), .CI(N2077));
ADDHX1 inst_cellmath__43_0_I1067 (.CO(N2258), .S(N3898), .A(N2966), .B(N3871));
ADDFXL inst_cellmath__43_0_I1068 (.CO(N3178), .S(N2714), .A(N3598), .B(N2680), .CI(N2398));
ADDFX1 inst_cellmath__43_0_I1069 (.CO(N4088), .S(N3641), .A(N2111), .B(N3301), .CI(N3014));
ADDFX1 inst_cellmath__43_0_I1070 (.CO(N2908), .S(N2453), .A(N2726), .B(N3919), .CI(N3642));
ADDFX1 inst_cellmath__43_0_I1071 (.CO(N3819), .S(N3366), .A(N3898), .B(N3334), .CI(N2154));
ADDFX1 inst_cellmath__43_0_I1072 (.CO(N2637), .S(N2188), .A(N2714), .B(N3065), .CI(N3978));
ADDFX1 inst_cellmath__43_0_I1073 (.CO(N3564), .S(N3102), .A(N2453), .B(N3641), .CI(N2790));
ADDFX1 inst_cellmath__43_0_I1074 (.CO(N2372), .S(N4010), .A(N3714), .B(N3366), .CI(N2188));
ADDFX1 inst_cellmath__43_0_I1075 (.CO(N3285), .S(N2825), .A(N2527), .B(N3102), .CI(N4010));
ADDHX1 inst_cellmath__43_0_I1076 (.CO(N2108), .S(N3745), .A(N3881), .B(N2689));
ADDFX1 inst_cellmath__43_0_I1077 (.CO(N3019), .S(N2559), .A(N2408), .B(N3606), .CI(N3311));
ADDFX1 inst_cellmath__43_0_I1078 (.CO(N3931), .S(N3483), .A(N2120), .B(N3025), .CI(N3929));
ADDFX1 inst_cellmath__43_0_I1079 (.CO(N2748), .S(N2294), .A(N2734), .B(N2455), .CI(N3652));
ADDFX1 inst_cellmath__43_0_I1080 (.CO(N3675), .S(N3210), .A(N2258), .B(N3360), .CI(N3745));
ADDFX1 inst_cellmath__43_0_I1081 (.CO(N2483), .S(N2029), .A(N4088), .B(N3178), .CI(N2908));
ADDFX1 inst_cellmath__43_0_I1082 (.CO(N3404), .S(N2943), .A(N3483), .B(N2559), .CI(N2294));
ADDFX1 inst_cellmath__43_0_I1083 (.CO(N2217), .S(N3851), .A(N3210), .B(N3819), .CI(N2029));
ADDFXL inst_cellmath__43_0_I1084 (.CO(N3130), .S(N2673), .A(N2637), .B(N3564), .CI(N2943));
ADDFX1 inst_cellmath__43_0_I1085 (.CO(N4048), .S(N3600), .A(N3851), .B(N2372), .CI(N2673));
ADDHX1 inst_cellmath__43_0_I1086 (.CO(N2866), .S(N2407), .A(N2698), .B(N3616));
ADDFX1 inst_cellmath__43_0_I1087 (.CO(N3776), .S(N3323), .A(N3321), .B(N2418), .CI(N2129));
ADDFX1 inst_cellmath__43_0_I1088 (.CO(N2599), .S(N2142), .A(N3938), .B(N3037), .CI(N2742));
ADDFX1 inst_cellmath__43_0_I1089 (.CO(N3519), .S(N3055), .A(N2465), .B(N3662), .CI(N3369));
ADDFX1 inst_cellmath__43_0_I1090 (.CO(N2330), .S(N3968), .A(N3085), .B(N2179), .CI(N2108));
ADDFX1 inst_cellmath__43_0_I1091 (.CO(N3246), .S(N2781), .A(N3019), .B(N2407), .CI(N3931));
ADDFX1 inst_cellmath__43_0_I1092 (.CO(N2068), .S(N3705), .A(N3323), .B(N2748), .CI(N2142));
ADDFX1 inst_cellmath__43_0_I1093 (.CO(N2973), .S(N2517), .A(N3675), .B(N3055), .CI(N2483));
ADDFX1 inst_cellmath__43_0_I1094 (.CO(N3890), .S(N3440), .A(N3404), .B(N3968), .CI(N2781));
ADDFX1 inst_cellmath__43_0_I1095 (.CO(N2707), .S(N2245), .A(N2517), .B(N3705), .CI(N2217));
ADDFX1 inst_cellmath__43_0_I1096 (.CO(N3634), .S(N3169), .A(N3130), .B(N3440), .CI(N2245));
ADDHX1 inst_cellmath__43_0_I1097 (.CO(N2445), .S(N4081), .A(N3627), .B(N2426));
ADDFXL inst_cellmath__43_0_I1098 (.CO(N3357), .S(N2896), .A(N3332), .B(N2140), .CI(N3043));
ADDFX1 inst_cellmath__43_0_I1099 (.CO(N2176), .S(N3811), .A(N3944), .B(N2751), .CI(N3671));
ADDFX1 inst_cellmath__43_0_I1100 (.CO(N3093), .S(N2629), .A(N3379), .B(N2473), .CI(N2189));
ADDFX1 inst_cellmath__43_0_I1101 (.CO(N4003), .S(N3551), .A(N3998), .B(N3094), .CI(N2800));
ADDFX1 inst_cellmath__43_0_I1102 (.CO(N2816), .S(N2362), .A(N4081), .B(N2866), .CI(N3776));
ADDFXL inst_cellmath__43_0_I1103 (.CO(N3737), .S(N3278), .A(N3519), .B(N2599), .CI(N2896));
ADDFXL inst_cellmath__43_0_I1104 (.CO(N2551), .S(N2097), .A(N3811), .B(N2330), .CI(N2629));
ADDFX1 inst_cellmath__43_0_I1105 (.CO(N3471), .S(N3009), .A(N3246), .B(N3551), .CI(N2068));
ADDFX1 inst_cellmath__43_0_I1106 (.CO(N2286), .S(N3921), .A(N3278), .B(N2362), .CI(N2097));
ADDFX1 inst_cellmath__43_0_I1107 (.CO(N3202), .S(N2738), .A(N3890), .B(N2973), .CI(N3009));
ADDFX1 inst_cellmath__43_0_I1108 (.CO(N2021), .S(N3667), .A(N2707), .B(N3921), .CI(N2738));
ADDHX1 inst_cellmath__43_0_I1109 (.CO(N2934), .S(N2474), .A(N2435), .B(N3340));
ADDFX1 inst_cellmath__43_0_I1110 (.CO(N3843), .S(N3394), .A(N3056), .B(N2152), .CI(N3952));
ADDFX1 inst_cellmath__43_0_I1111 (.CO(N2663), .S(N2209), .A(N3678), .B(N2759), .CI(N2480));
ADDFX1 inst_cellmath__43_0_I1112 (.CO(N3591), .S(N3122), .A(N2197), .B(N3388), .CI(N3104));
ADDFX1 inst_cellmath__43_0_I1113 (.CO(N2397), .S(N4035), .A(N2810), .B(N4005), .CI(N3721));
ADDFX1 inst_cellmath__43_0_I1114 (.CO(N3313), .S(N2852), .A(N2445), .B(N2528), .CI(N2474));
ADDFXL inst_cellmath__43_0_I1115 (.CO(N2131), .S(N3765), .A(N3093), .B(N3357), .CI(N2176));
ADDFX1 inst_cellmath__43_0_I1116 (.CO(N3042), .S(N2588), .A(N3394), .B(N4003), .CI(N2209));
ADDFX1 inst_cellmath__43_0_I1117 (.CO(N3955), .S(N3507), .A(N4035), .B(N3122), .CI(N2816));
ADDFX1 inst_cellmath__43_0_I1118 (.CO(N2768), .S(N2318), .A(N2852), .B(N3737), .CI(N3765));
ADDFX1 inst_cellmath__43_0_I1119 (.CO(N3693), .S(N3235), .A(N2588), .B(N2551), .CI(N3471));
ADDFX1 inst_cellmath__43_0_I1120 (.CO(N2508), .S(N2057), .A(N2286), .B(N3507), .CI(N2318));
ADDFX1 inst_cellmath__43_0_I1121 (.CO(N3429), .S(N2963), .A(N3235), .B(N3202), .CI(N2057));
ADDHX1 inst_cellmath__43_0_I1122 (.CO(N2236), .S(N3880), .A(N3351), .B(N2163));
ADDFXL inst_cellmath__43_0_I1123 (.CO(N3159), .S(N2696), .A(N3066), .B(N3965), .CI(N2766));
ADDFX1 inst_cellmath__43_0_I1124 (.CO(N4071), .S(N3624), .A(N2488), .B(N3687), .CI(N3398));
ADDFX1 inst_cellmath__43_0_I1125 (.CO(N2886), .S(N2434), .A(N3113), .B(N2205), .CI(N4014));
ADDFX1 inst_cellmath__43_0_I1126 (.CO(N3802), .S(N3350), .A(N3730), .B(N2819), .CI(N2537));
ADDFX1 inst_cellmath__43_0_I1127 (.CO(N2620), .S(N2168), .A(N2246), .B(N3448), .CI(N2934));
ADDFX1 inst_cellmath__43_0_I1128 (.CO(N3542), .S(N3084), .A(N3843), .B(N3880), .CI(N2663));
ADDFXL inst_cellmath__43_0_I1129 (.CO(N2354), .S(N3994), .A(N2397), .B(N3591), .CI(N2696));
ADDFX1 inst_cellmath__43_0_I1130 (.CO(N3270), .S(N2807), .A(N2434), .B(N3624), .CI(N3350));
ADDFX1 inst_cellmath__43_0_I1131 (.CO(N2087), .S(N3729), .A(N2168), .B(N3313), .CI(N2131));
ADDFX1 inst_cellmath__43_0_I1132 (.CO(N3002), .S(N2544), .A(N3084), .B(N3042), .CI(N3994));
ADDFX1 inst_cellmath__43_0_I1133 (.CO(N3912), .S(N3461), .A(N3955), .B(N2807), .CI(N3729));
ADDFX1 inst_cellmath__43_0_I1134 (.CO(N2728), .S(N2276), .A(N2544), .B(N2768), .CI(N3693));
ADDFX1 inst_cellmath__43_0_I1135 (.CO(N3657), .S(N3196), .A(N2508), .B(N3461), .CI(N2276));
ADDHX1 inst_cellmath__43_0_I1136 (.CO(N2468), .S(N2011), .A(N2171), .B(N3076));
ADDFX1 inst_cellmath__43_0_I1137 (.CO(N3382), .S(N2925), .A(N2779), .B(N3976), .CI(N3695));
ADDFX1 inst_cellmath__43_0_I1138 (.CO(N2202), .S(N3836), .A(N3409), .B(N2499), .CI(N2213));
ADDFX1 inst_cellmath__43_0_I1139 (.CO(N3116), .S(N2652), .A(N4021), .B(N3121), .CI(N2826));
ADDFX1 inst_cellmath__43_0_I1140 (.CO(N4026), .S(N3582), .A(N2547), .B(N3738), .CI(N3456));
ADDFX1 inst_cellmath__43_0_I1141 (.CO(N2841), .S(N2389), .A(N3166), .B(N2255), .CI(N4072));
ADDFX1 inst_cellmath__43_0_I1142 (.CO(N3757), .S(N3303), .A(N2011), .B(N2236), .CI(N3159));
ADDFX1 inst_cellmath__43_0_I1143 (.CO(N2577), .S(N2122), .A(N2886), .B(N4071), .CI(N3802));
ADDFX1 inst_cellmath__43_0_I1144 (.CO(N3498), .S(N3036), .A(N3836), .B(N2925), .CI(N2620));
ADDFX1 inst_cellmath__43_0_I1145 (.CO(N2310), .S(N3946), .A(N3582), .B(N2652), .CI(N2389));
ADDFX1 inst_cellmath__43_0_I1146 (.CO(N3228), .S(N2761), .A(N2354), .B(N3542), .CI(N3270));
ADDFX1 inst_cellmath__43_0_I1147 (.CO(N2046), .S(N3686), .A(N3303), .B(N2122), .CI(N3036));
ADDFX1 inst_cellmath__43_0_I1148 (.CO(N2956), .S(N2501), .A(N2087), .B(N3946), .CI(N3002));
ADDFX1 inst_cellmath__43_0_I1149 (.CO(N3869), .S(N3420), .A(N3686), .B(N2761), .CI(N3912));
ADDFX1 inst_cellmath__43_0_I1150 (.CO(N2688), .S(N2230), .A(N2728), .B(N2501), .CI(N3420));
ADDHX1 inst_cellmath__43_0_I1151 (.CO(N3613), .S(N3148), .A(N3086), .B(N3986));
ADDFXL inst_cellmath__43_0_I1152 (.CO(N2424), .S(N4065), .A(N3706), .B(N2791), .CI(N2506));
ADDFXL inst_cellmath__43_0_I1153 (.CO(N3339), .S(N2879), .A(N2224), .B(N3418), .CI(N3128));
ADDFX1 inst_cellmath__43_0_I1154 (.CO(N2160), .S(N3793), .A(N2837), .B(N4030), .CI(N3747));
ADDFX1 inst_cellmath__43_0_I1155 (.CO(N3074), .S(N2611), .A(N3463), .B(N2554), .CI(N2265));
ADDFX1 inst_cellmath__43_0_I1156 (.CO(N3985), .S(N3533), .A(N4082), .B(N3179), .CI(N2887));
ADDFX1 inst_cellmath__43_0_I1157 (.CO(N2796), .S(N2346), .A(N2468), .B(N3790), .CI(N3148));
ADDFX1 inst_cellmath__43_0_I1158 (.CO(N3720), .S(N3261), .A(N2202), .B(N3382), .CI(N3116));
ADDFXL inst_cellmath__43_0_I1159 (.CO(N2532), .S(N2079), .A(N2841), .B(N4026), .CI(N4065));
ADDFX1 inst_cellmath__43_0_I1160 (.CO(N3453), .S(N2994), .A(N3793), .B(N2879), .CI(N2611));
ADDFX1 inst_cellmath__43_0_I1161 (.CO(N2264), .S(N3903), .A(N2577), .B(N3533), .CI(N3757));
ADDFX1 inst_cellmath__43_0_I1162 (.CO(N3186), .S(N2719), .A(N3498), .B(N2346), .CI(N3261));
ADDFX1 inst_cellmath__43_0_I1163 (.CO(N4096), .S(N3647), .A(N2079), .B(N2310), .CI(N2994));
ADDFX1 inst_cellmath__43_0_I1164 (.CO(N2913), .S(N2460), .A(N3903), .B(N3228), .CI(N2046));
ADDFX1 inst_cellmath__43_0_I1165 (.CO(N3827), .S(N3372), .A(N3647), .B(N2719), .CI(N2956));
ADDFX1 inst_cellmath__43_0_I1166 (.CO(N2644), .S(N2194), .A(N3869), .B(N2460), .CI(N3372));
ADDHX1 inst_cellmath__43_0_I1167 (.CO(N3570), .S(N3107), .A(N3996), .B(N2801));
ADDFX1 inst_cellmath__43_0_I1168 (.CO(N2380), .S(N4016), .A(N2515), .B(N3715), .CI(N3427));
ADDFX1 inst_cellmath__43_0_I1169 (.CO(N3291), .S(N2832), .A(N3136), .B(N2231), .CI(N4040));
ADDFX1 inst_cellmath__43_0_I1170 (.CO(N2114), .S(N3750), .A(N2846), .B(N2563), .CI(N3756));
ADDFX1 inst_cellmath__43_0_I1171 (.CO(N3028), .S(N2566), .A(N2278), .B(N3472), .CI(N3190));
ADDFX1 inst_cellmath__43_0_I1172 (.CO(N3937), .S(N3490), .A(N2897), .B(N4089), .CI(N3799));
ADDFX1 inst_cellmath__43_0_I1173 (.CO(N2754), .S(N2300), .A(N3524), .B(N2612), .CI(N3613));
ADDFX1 inst_cellmath__43_0_I1174 (.CO(N3681), .S(N3215), .A(N3107), .B(N3339), .CI(N2424));
ADDFX1 inst_cellmath__43_0_I1175 (.CO(N2487), .S(N2037), .A(N3074), .B(N2160), .CI(N3985));
ADDFX1 inst_cellmath__43_0_I1176 (.CO(N3412), .S(N2949), .A(N2832), .B(N4016), .CI(N3750));
ADDFX1 inst_cellmath__43_0_I1177 (.CO(N2223), .S(N3857), .A(N3490), .B(N2566), .CI(N2796));
ADDFX1 inst_cellmath__43_0_I1178 (.CO(N3140), .S(N2678), .A(N3720), .B(N2300), .CI(N2532));
ADDFX1 inst_cellmath__43_0_I1179 (.CO(N4054), .S(N3605), .A(N2037), .B(N3453), .CI(N3215));
ADDFX1 inst_cellmath__43_0_I1180 (.CO(N2871), .S(N2416), .A(N2264), .B(N2949), .CI(N3857));
ADDFX1 inst_cellmath__43_0_I1181 (.CO(N3785), .S(N3331), .A(N2678), .B(N3186), .CI(N4096));
ADDFX1 inst_cellmath__43_0_I1182 (.CO(N2605), .S(N2149), .A(N2416), .B(N3605), .CI(N2913));
ADDFX1 inst_cellmath__43_0_I1183 (.CO(N3523), .S(N3064), .A(N3827), .B(N3331), .CI(N2149));
ADDHX1 inst_cellmath__43_0_I1184 (.CO(N2338), .S(N3975), .A(N2811), .B(N3722));
ADDFXL inst_cellmath__43_0_I1185 (.CO(N3252), .S(N2787), .A(N3438), .B(N2524), .CI(N2237));
ADDFX1 inst_cellmath__43_0_I1186 (.CO(N2071), .S(N3713), .A(N4051), .B(N3146), .CI(N2860));
ADDFX1 inst_cellmath__43_0_I1187 (.CO(N2983), .S(N2523), .A(N2573), .B(N3764), .CI(N3485));
ADDFX1 inst_cellmath__43_0_I1188 (.CO(N3895), .S(N3445), .A(N4100), .B(N2287), .CI(N3198));
ADDFXL inst_cellmath__43_0_I1189 (.CO(N2710), .S(N2254), .A(N2905), .B(N2621), .CI(N3808));
ADDFX1 inst_cellmath__43_0_I1190 (.CO(N3639), .S(N3174), .A(N3240), .B(N2334), .CI(N3534));
ADDFX1 inst_cellmath__43_0_I1191 (.CO(N2449), .S(N4085), .A(N3975), .B(N3570), .CI(N2380));
ADDFX1 inst_cellmath__43_0_I1192 (.CO(N3363), .S(N2904), .A(N2114), .B(N3028), .CI(N3291));
ADDFX1 inst_cellmath__43_0_I1193 (.CO(N2185), .S(N3816), .A(N2787), .B(N3937), .CI(N2754));
ADDFX1 inst_cellmath__43_0_I1194 (.CO(N3098), .S(N2634), .A(N2523), .B(N3713), .CI(N3445));
ADDFXL inst_cellmath__43_0_I1195 (.CO(N4006), .S(N3560), .A(N2254), .B(N3174), .CI(N3681));
ADDFX1 inst_cellmath__43_0_I1196 (.CO(N2823), .S(N2370), .A(N3412), .B(N2487), .CI(N4085));
ADDFX1 inst_cellmath__43_0_I1197 (.CO(N3742), .S(N3282), .A(N2223), .B(N2904), .CI(N3816));
ADDFX1 inst_cellmath__43_0_I1198 (.CO(N2555), .S(N2104), .A(N2634), .B(N3140), .CI(N3560));
ADDFX1 inst_cellmath__43_0_I1199 (.CO(N3478), .S(N3016), .A(N2370), .B(N4054), .CI(N2871));
ADDFX1 inst_cellmath__43_0_I1200 (.CO(N2290), .S(N3928), .A(N3282), .B(N2104), .CI(N3785));
ADDFX1 inst_cellmath__43_0_I1201 (.CO(N3207), .S(N2745), .A(N2605), .B(N3016), .CI(N3928));
ADDHXL inst_cellmath__43_0_I1202 (.CO(N2026), .S(N3673), .A(N3731), .B(N2534));
ADDFXL inst_cellmath__43_0_I1203 (.CO(N2938), .S(N2479), .A(N2247), .B(N3449), .CI(N3156));
ADDFXL inst_cellmath__43_0_I1204 (.CO(N3848), .S(N3400), .A(N2872), .B(N4063), .CI(N3774));
ADDFXL inst_cellmath__43_0_I1205 (.CO(N2670), .S(N2215), .A(N3494), .B(N2582), .CI(N2296));
ADDFX1 inst_cellmath__43_0_I1206 (.CO(N3596), .S(N3127), .A(N2914), .B(N3206), .CI(N2013));
ADDFX1 inst_cellmath__43_0_I1207 (.CO(N2404), .S(N4043), .A(N2630), .B(N3820), .CI(N3543));
ADDFX1 inst_cellmath__43_0_I1208 (.CO(N3320), .S(N2863), .A(N2343), .B(N3253), .CI(N2065));
ADDFX1 inst_cellmath__43_0_I1209 (.CO(N2139), .S(N3773), .A(N2338), .B(N2961), .CI(N3673));
ADDFHXL inst_cellmath__43_0_I1210 (.CO(N3052), .S(N2596), .A(N2983), .B(N3252), .CI(N2071));
ADDFX1 inst_cellmath__43_0_I1211 (.CO(N3962), .S(N3517), .A(N2710), .B(N3895), .CI(N3639));
ADDFXL inst_cellmath__43_0_I1212 (.CO(N2778), .S(N2326), .A(N2215), .B(N2479), .CI(N3400));
ADDFX1 inst_cellmath__43_0_I1213 (.CO(N3702), .S(N3244), .A(N4043), .B(N3127), .CI(N2863));
ADDFX1 inst_cellmath__43_0_I1214 (.CO(N2514), .S(N2064), .A(N2449), .B(N3363), .CI(N3773));
ADDFHX1 inst_cellmath__43_0_I1215 (.CO(N3436), .S(N2969), .A(N2596), .B(N2185), .CI(N3517));
ADDFX1 inst_cellmath__43_0_I1216 (.CO(N2244), .S(N3887), .A(N4006), .B(N3098), .CI(N2326));
ADDFX1 inst_cellmath__43_0_I1217 (.CO(N3165), .S(N2703), .A(N2064), .B(N3244), .CI(N2823));
ADDFX1 inst_cellmath__43_0_I1218 (.CO(N4078), .S(N3633), .A(N2969), .B(N3742), .CI(N2555));
ADDFX1 inst_cellmath__43_0_I1219 (.CO(N2894), .S(N2440), .A(N3478), .B(N3887), .CI(N2703));
ADDFXL inst_cellmath__43_0_I1220 (.CO(N3807), .S(N3354), .A(N2290), .B(N3633), .CI(N2440));
ADDHX1 inst_cellmath__43_0_I1221 (.CO(N2627), .S(N2175), .A(N2545), .B(N3457));
ADDFHXL inst_cellmath__43_0_I1222 (.CO(N3550), .S(N3090), .A(N2256), .B(N3167), .CI(N4069));
ADDFHX1 inst_cellmath__43_0_I1223 (.CO(N2359), .S(N4000), .A(N3781), .B(N2880), .CI(N2593));
ADDFXL inst_cellmath__43_0_I1224 (.CO(N3276), .S(N2815), .A(N2308), .B(N3213), .CI(N3503));
ADDFXL inst_cellmath__43_0_I1225 (.CO(N2094), .S(N3734), .A(N2926), .B(N2022), .CI(N3830));
ADDFX1 inst_cellmath__43_0_I1226 (.CO(N3007), .S(N2549), .A(N2351), .B(N3552), .CI(N2638));
ADDFX1 inst_cellmath__43_0_I1227 (.CO(N3918), .S(N3469), .A(N2072), .B(N3262), .CI(N2970));
ADDFXL inst_cellmath__43_0_I1228 (.CO(N2735), .S(N2283), .A(N2686), .B(N3873), .CI(N2026));
ADDFX1 inst_cellmath__43_0_I1229 (.CO(N3664), .S(N3200), .A(N2175), .B(N2938), .CI(N3848));
ADDFXL inst_cellmath__43_0_I1230 (.CO(N2472), .S(N2018), .A(N2670), .B(N3596), .CI(N2404));
ADDFXL inst_cellmath__43_0_I1231 (.CO(N3390), .S(N2929), .A(N3090), .B(N3320), .CI(N4000));
ADDFHXL inst_cellmath__43_0_I1232 (.CO(N2206), .S(N3841), .A(N2815), .B(N3734), .CI(N2549));
ADDFX1 inst_cellmath__43_0_I1233 (.CO(N3120), .S(N2660), .A(N2139), .B(N3469), .CI(N3052));
ADDFHXL inst_cellmath__43_0_I1234 (.CO(N4032), .S(N3586), .A(N3962), .B(N2283), .CI(N2778));
ADDFX1 inst_cellmath__43_0_I1235 (.CO(N2848), .S(N2395), .A(N2018), .B(N3702), .CI(N3200));
ADDFXL inst_cellmath__43_0_I1236 (.CO(N3763), .S(N3310), .A(N3841), .B(N2929), .CI(N2514));
ADDFHXL inst_cellmath__43_0_I1237 (.CO(N2584), .S(N2127), .A(N2660), .B(N3436), .CI(N3586));
ADDFXL inst_cellmath__43_0_I1238 (.CO(N3504), .S(N3041), .A(N2395), .B(N2244), .CI(N3310));
ADDFX1 inst_cellmath__43_0_I1239 (.CO(N2315), .S(N3951), .A(N2127), .B(N3165), .CI(N4078));
ADDFHXL inst_cellmath__43_0_I1240 (.CO(N3233), .S(N2764), .A(N2894), .B(N3041), .CI(N3951));
XNOR2X1 inst_cellmath__43_0_I1241 (.Y(N3692), .A(N3464), .B(N2266));
OR2XL inst_cellmath__43_0_I1242 (.Y(N2053), .A(N2266), .B(N3464));
ADDFXL inst_cellmath__43_0_I1243 (.CO(N3877), .S(N3425), .A(N4079), .B(N3176), .CI(N2888));
ADDFHXL inst_cellmath__43_0_I1244 (.CO(N2692), .S(N2235), .A(N2602), .B(N3514), .CI(N3791));
ADDFHXL inst_cellmath__43_0_I1245 (.CO(N3619), .S(N3155), .A(N2316), .B(N2030), .CI(N3224));
ADDFXL inst_cellmath__43_0_I1246 (.CO(N2432), .S(N4067), .A(N3839), .B(N2935), .CI(N2648));
ADDFHXL inst_cellmath__43_0_I1247 (.CO(N3345), .S(N2885), .A(N2363), .B(N3561), .CI(N3271));
ADDFXL inst_cellmath__43_0_I1248 (.CO(N2165), .S(N3798), .A(N2979), .B(N2080), .CI(N3888));
ADDFX1 inst_cellmath__43_0_I1249 (.CO(N3082), .S(N2616), .A(N2410), .B(N3611), .CI(N2693));
ADDFHXL inst_cellmath__43_0_I1250 (.CO(N3990), .S(N3539), .A(N3692), .B(N2627), .CI(N3550));
ADDFHXL inst_cellmath__43_0_I1251 (.CO(N2804), .S(N2350), .A(N2094), .B(N2359), .CI(N3276));
ADDFXL inst_cellmath__43_0_I1252 (.CO(N3726), .S(N3266), .A(N3918), .B(N3007), .CI(N3425));
ADDFX1 inst_cellmath__43_0_I1253 (.CO(N2539), .S(N2086), .A(N3155), .B(N2235), .CI(N2735));
ADDFX1 inst_cellmath__43_0_I1254 (.CO(N3460), .S(N2998), .A(N2885), .B(N4067), .CI(N3798));
ADDFX1 inst_cellmath__43_0_I1255 (.CO(N2272), .S(N3908), .A(N3664), .B(N2616), .CI(N2472));
ADDFXL inst_cellmath__43_0_I1256 (.CO(N3191), .S(N2727), .A(N2350), .B(N3539), .CI(N3390));
ADDFX1 inst_cellmath__43_0_I1257 (.CO(N4105), .S(N3653), .A(N3266), .B(N2206), .CI(N2086));
ADDFX1 inst_cellmath__43_0_I1258 (.CO(N2919), .S(N2464), .A(N2998), .B(N3120), .CI(N4032));
ADDFXL inst_cellmath__43_0_I1259 (.CO(N3831), .S(N3381), .A(N2848), .B(N3908), .CI(N2727));
ADDFXL inst_cellmath__43_0_I1261 (.CO(N3577), .S(N3112), .A(N3381), .B(N2464), .CI(N3504));
ADDFHXL inst_cellmath__43_0_I11173 (.CO(N18827), .S(N2198), .A(N3653), .B(N3763), .CI(N2584));
ADDFXL inst_cellmath__43_0_I1262 (.CO(N2385), .S(N4022), .A(N2315), .B(N2198), .CI(N3112));
ADDHXL inst_cellmath__43_0_I1263 (.CO(N3299), .S(N2838), .A(N2400), .B(N3187));
ADDFXL inst_cellmath__43_0_I1264 (.CO(N2118), .S(N3755), .A(N4090), .B(N2279), .CI(N2898));
ADDFX1 inst_cellmath__43_0_I1265 (.CO(N3034), .S(N2574), .A(N2609), .B(N3800), .CI(N3525));
ADDFHXL inst_cellmath__43_0_I1266 (.CO(N3943), .S(N3495), .A(N3231), .B(N2042), .CI(N2327));
ADDFX1 inst_cellmath__43_0_I1267 (.CO(N2758), .S(N2306), .A(N3847), .B(N2655), .CI(N2946));
ADDFX1 inst_cellmath__43_0_I1268 (.CO(N3685), .S(N3225), .A(N2373), .B(N3572), .CI(N3279));
ADDFX1 inst_cellmath__43_0_I1269 (.CO(N2497), .S(N2043), .A(N2991), .B(N2088), .CI(N3896));
ADDFX1 inst_cellmath__43_0_I1270 (.CO(N3416), .S(N2954), .A(N3620), .B(N2704), .CI(N2420));
ADDFXL inst_cellmath__43_0_I1271 (.CO(N2229), .S(N3867), .A(N2053), .B(N3327), .CI(N2838));
ADDFHXL inst_cellmath__43_0_I1272 (.CO(N3145), .S(N2685), .A(N3619), .B(N2692), .CI(N3877));
ADDFXL inst_cellmath__43_0_I1273 (.CO(N4061), .S(N3610), .A(N3345), .B(N2432), .CI(N2165));
ADDFX1 inst_cellmath__43_0_I1274 (.CO(N2877), .S(N2422), .A(N3082), .B(N3755), .CI(N2574));
ADDFX1 inst_cellmath__43_0_I1275 (.CO(N3789), .S(N3336), .A(N3225), .B(N3495), .CI(N2306));
ADDFXL inst_cellmath__43_0_I1276 (.CO(N2608), .S(N2157), .A(N2954), .B(N2043), .CI(N3990));
ADDFX1 inst_cellmath__43_0_I1277 (.CO(N3532), .S(N3071), .A(N2804), .B(N3867), .CI(N3726));
ADDFXL inst_cellmath__43_0_I1278 (.CO(N2341), .S(N3982), .A(N2539), .B(N2685), .CI(N3610));
ADDFXL inst_cellmath__43_0_I1279 (.CO(N3258), .S(N2794), .A(N2422), .B(N3460), .CI(N3336));
ADDFXL inst_cellmath__43_0_I11176 (.CO(N18841), .S(N3451), .A(N2919), .B(N2794), .CI(N3831));
ADDFX1 inst_cellmath__43_0_I11175 (.CO(N18820), .S(N18857), .A(N4105), .B(N3071), .CI(N3982));
ADDFX1 inst_cellmath__43_0_I11174 (.CO(N18848), .S(N18836), .A(N2157), .B(N2272), .CI(N3191));
ADDFHXL inst_cellmath__43_0_I11177 (.CO(N18814), .S(N2260), .A(N18857), .B(N18836), .CI(N18827));
ADDFHX1 inst_cellmath__43_0_I1284 (.CO(N3643), .S(N3182), .A(N3577), .B(N3451), .CI(N2260));
ADDHX1 inst_cellmath__43_0_I1285 (.CO(N2456), .S(N4093), .A(N3317), .B(N2906));
ADDFHXL inst_cellmath__43_0_I1286 (.CO(N3368), .S(N2910), .A(N4101), .B(N3809), .CI(N2618));
ADDFHXL inst_cellmath__43_0_I1287 (.CO(N2190), .S(N3823), .A(N2335), .B(N3535), .CI(N3241));
ADDFHX1 inst_cellmath__43_0_I1288 (.CO(N3103), .S(N2641), .A(N3854), .B(N2955), .CI(N2052));
ADDFHXL inst_cellmath__43_0_I1289 (.CO(N4013), .S(N3566), .A(N2664), .B(N3583), .CI(N2383));
ADDFXL inst_cellmath__43_0_I1290 (.CO(N2827), .S(N2374), .A(N3000), .B(N2095), .CI(N3286));
ADDFXL inst_cellmath__43_0_I1291 (.CO(N3746), .S(N3289), .A(N2711), .B(N3904), .CI(N3630));
ADDFX1 inst_cellmath__43_0_I1292 (.CO(N2564), .S(N2109), .A(N2146), .B(N2429), .CI(N3337));
ADDFXL inst_cellmath__43_0_I1293 (.CO(N3486), .S(N3022), .A(N4093), .B(N3299), .CI(N2118));
ADDFHXL inst_cellmath__43_0_I1294 (.CO(N2295), .S(N3935), .A(N2758), .B(N3034), .CI(N3943));
ADDFHXL inst_cellmath__43_0_I1295 (.CO(N3214), .S(N2749), .A(N2497), .B(N3685), .CI(N3416));
ADDFX1 inst_cellmath__43_0_I1296 (.CO(N2032), .S(N3677), .A(N2641), .B(N3823), .CI(N2910));
ADDFX1 inst_cellmath__43_0_I1297 (.CO(N2945), .S(N2486), .A(N3566), .B(N2374), .CI(N3289));
ADDFXL inst_cellmath__43_0_I1298 (.CO(N3855), .S(N3407), .A(N2229), .B(N2109), .CI(N3145));
ADDFX1 inst_cellmath__43_0_I1299 (.CO(N2675), .S(N2220), .A(N3022), .B(N4061), .CI(N3935));
ADDFXL inst_cellmath__43_0_I1300 (.CO(N3601), .S(N3134), .A(N2877), .B(N2749), .CI(N3789));
ADDFXL inst_cellmath__43_0_I1307 (.CO(N3711), .S(N3249), .A(N3817), .B(N2134), .CI(N2631));
ADDFHXL inst_cellmath__43_0_I1308 (.CO(N2520), .S(N2070), .A(N2344), .B(N3544), .CI(N3250));
ADDFXL inst_cellmath__43_0_I1309 (.CO(N3443), .S(N2978), .A(N2962), .B(N3866), .CI(N2066));
ADDFXL inst_cellmath__43_0_I1310 (.CO(N2250), .S(N3892), .A(N3594), .B(N2674), .CI(N2393));
ADDFXL inst_cellmath__43_0_I1311 (.CO(N3171), .S(N2709), .A(N2105), .B(N3295), .CI(N3010));
ADDFXL inst_cellmath__43_0_I1312 (.CO(N4083), .S(N3636), .A(N2720), .B(N3913), .CI(N3637));
ADDFX1 inst_cellmath__43_0_I1313 (.CO(N2902), .S(N2447), .A(N3346), .B(N2441), .CI(N2158));
ADDFHXL inst_cellmath__43_0_I1314 (.CO(N3813), .S(N3359), .A(N2456), .B(N3058), .CI(N3368));
ADDFHXL inst_cellmath__43_0_I1315 (.CO(N2632), .S(N2181), .A(N3103), .B(N4013), .CI(N2190));
ADDFXL inst_cellmath__43_0_I1316 (.CO(N3557), .S(N3096), .A(N2564), .B(N2827), .CI(N3746));
ADDFXL inst_cellmath__43_0_I1317 (.CO(N2365), .S(N4004), .A(N3249), .B(N2070), .CI(N2978));
ADDFX1 inst_cellmath__43_0_I1318 (.CO(N3280), .S(N2820), .A(N3636), .B(N3892), .CI(N2709));
ADDFHXL inst_cellmath__43_0_I1319 (.CO(N2101), .S(N3740), .A(N3486), .B(N2447), .CI(N2295));
ADDFHXL inst_cellmath__43_0_I1320 (.CO(N3011), .S(N2553), .A(N3214), .B(N3359), .CI(N2032));
ADDFXL inst_cellmath__43_0_I1321 (.CO(N3925), .S(N3473), .A(N2181), .B(N2945), .CI(N3096));
ADDFX1 inst_cellmath__43_0_I1322 (.CO(N2741), .S(N2288), .A(N2820), .B(N3855), .CI(N4004));
ADDFHXL inst_cellmath__43_0_I1323 (.CO(N3669), .S(N3205), .A(N3740), .B(N2675), .CI(N3601));
ADDFX1 inst_cellmath__43_0_I11178 (.CO(N2412), .S(N18825), .A(N3677), .B(N2486), .CI(N2608));
ADDFHXL inst_cellmath__43_0_I1324 (.CO(N2477), .S(N2023), .A(N3473), .B(N2553), .CI(N2412));
ADDFHXL inst_cellmath__43_0_I11179 (.CO(N3326), .S(N18846), .A(N3532), .B(N3407), .CI(N2341));
ADDFHXL inst_cellmath__43_0_I1325 (.CO(N3396), .S(N2936), .A(N3326), .B(N2288), .CI(N3205));
ADDFXL inst_cellmath__43_0_I11180 (.CO(N2145), .S(N18818), .A(N3134), .B(N2220), .CI(N3258));
ADDFHXL inst_cellmath__43_0_I11181 (.CO(N3060), .S(N18839), .A(N18848), .B(N18825), .CI(N18846));
ADDFHXL inst_cellmath__43_0_I1326 (.CO(N2212), .S(N3846), .A(N2023), .B(N2145), .CI(N3060));
ADDFHXL inst_cellmath__43_0_I11182 (.CO(N18823), .S(N18860), .A(N18818), .B(N18820), .CI(N18841));
ADDFHXL inst_cellmath__43_0_I11183 (.CO(N2783), .S(N2333), .A(N18814), .B(N18839), .CI(N18860));
ADDFHXL inst_cellmath__43_0_I11184 (.CO(N3125), .S(N2666), .A(N18823), .B(N2936), .CI(N3846));
NAND2X2 inst_cellmath__43_0_I11185 (.Y(N2701), .A(N2783), .B(N2666));
INVXL buf1_A_I4232 (.Y(N9406), .A(N2666));
INVX1 buf1_A_I4233 (.Y(N3048), .A(N9406));
ADDFHXL inst_cellmath__43_0_I1330 (.CO(N4039), .S(N3593), .A(N3553), .B(N3046), .CI(N2352));
ADDFXL inst_cellmath__43_0_I1331 (.CO(N2856), .S(N2403), .A(N2073), .B(N3259), .CI(N2971));
ADDFXL inst_cellmath__43_0_I1332 (.CO(N3771), .S(N3316), .A(N2684), .B(N3874), .CI(N3602));
ADDFX1 inst_cellmath__43_0_I1333 (.CO(N2591), .S(N2133), .A(N3304), .B(N2401), .CI(N2115));
ADDFXL inst_cellmath__43_0_I1334 (.CO(N3512), .S(N3050), .A(N3922), .B(N3020), .CI(N2729));
ADDFXL inst_cellmath__43_0_I1335 (.CO(N2325), .S(N3958), .A(N2450), .B(N3644), .CI(N3355));
ADDFX1 inst_cellmath__43_0_I1336 (.CO(N3238), .S(N2770), .A(N3069), .B(N2166), .CI(N3972));
ADDFXL inst_cellmath__43_0_I1337 (.CO(N2060), .S(N3701), .A(N3711), .B(N2520), .CI(N3443));
ADDFXL inst_cellmath__43_0_I1338 (.CO(N2968), .S(N2511), .A(N4083), .B(N3171), .CI(N2250));
ADDFX1 inst_cellmath__43_0_I1339 (.CO(N3883), .S(N3430), .A(N2902), .B(N3593), .CI(N2403));
ADDFX1 inst_cellmath__43_0_I1340 (.CO(N2699), .S(N2241), .A(N3316), .B(N3050), .CI(N2133));
ADDFXL inst_cellmath__43_0_I1341 (.CO(N3629), .S(N3161), .A(N2770), .B(N3958), .CI(N3813));
ADDFX1 inst_cellmath__43_0_I1342 (.CO(N2437), .S(N4074), .A(N3557), .B(N2632), .CI(N2365));
ADDFX1 inst_cellmath__43_0_I1343 (.CO(N3352), .S(N2892), .A(N3280), .B(N2511), .CI(N3701));
ADDFX1 inst_cellmath__43_0_I1344 (.CO(N2173), .S(N3804), .A(N3430), .B(N2101), .CI(N2241));
ADDFXL inst_cellmath__43_0_I1345 (.CO(N3088), .S(N2622), .A(N3161), .B(N3011), .CI(N3925));
ADDFXL inst_cellmath__43_0_I1346 (.CO(N3997), .S(N3549), .A(N4074), .B(N2892), .CI(N2741));
ADDFXL inst_cellmath__43_0_I1347 (.CO(N2813), .S(N2356), .A(N3804), .B(N3669), .CI(N2622));
ADDFHXL inst_cellmath__43_0_I1348 (.CO(N3733), .S(N3273), .A(N3549), .B(N2477), .CI(N3396));
ADDFHX1 inst_cellmath__43_0_I1349 (.CO(N2546), .S(N2092), .A(N2212), .B(N2356), .CI(N3273));
ADDFX1 inst_cellmath__43_0_I1350 (.CO(N3467), .S(N3004), .A(N3959), .B(N2081), .CI(N3268));
ADDFXL inst_cellmath__43_0_I1351 (.CO(N2281), .S(N3914), .A(N2980), .B(N2691), .CI(N3885));
ADDFX1 inst_cellmath__43_0_I1352 (.CO(N3197), .S(N2733), .A(N2411), .B(N3612), .CI(N3314));
ADDFX1 inst_cellmath__43_0_I1353 (.CO(N2015), .S(N3660), .A(N3032), .B(N2123), .CI(N3932));
ADDFX1 inst_cellmath__43_0_I1354 (.CO(N2928), .S(N2470), .A(N3655), .B(N2736), .CI(N2461));
ADDFX1 inst_cellmath__43_0_I1355 (.CO(N3838), .S(N3387), .A(N2174), .B(N3364), .CI(N3080));
ADDFXL inst_cellmath__43_0_I1356 (.CO(N2657), .S(N2204), .A(N2784), .B(N3983), .CI(N4039));
ADDFXL inst_cellmath__43_0_I1357 (.CO(N3585), .S(N3118), .A(N3771), .B(N2856), .CI(N2591));
ADDFX1 inst_cellmath__43_0_I1358 (.CO(N2392), .S(N4029), .A(N2325), .B(N3512), .CI(N3238));
ADDFXL inst_cellmath__43_0_I1359 (.CO(N3307), .S(N2845), .A(N2733), .B(N3914), .CI(N3004));
ADDFX1 inst_cellmath__43_0_I1360 (.CO(N2125), .S(N3761), .A(N2470), .B(N3660), .CI(N3387));
ADDFX1 inst_cellmath__43_0_I1361 (.CO(N3039), .S(N2580), .A(N2968), .B(N2060), .CI(N2204));
ADDFHXL inst_cellmath__43_0_I1362 (.CO(N3949), .S(N3502), .A(N2699), .B(N3883), .CI(N3118));
ADDFX1 inst_cellmath__43_0_I1363 (.CO(N2763), .S(N2314), .A(N3629), .B(N4029), .CI(N2845));
ADDFHXL inst_cellmath__43_0_I1364 (.CO(N3689), .S(N3230), .A(N2437), .B(N3761), .CI(N3352));
ADDFHXL inst_cellmath__43_0_I1365 (.CO(N2504), .S(N2050), .A(N3502), .B(N2580), .CI(N2173));
ADDFHXL inst_cellmath__43_0_I1366 (.CO(N3422), .S(N2958), .A(N3088), .B(N2314), .CI(N3230));
ADDFHXL inst_cellmath__43_0_I1367 (.CO(N2233), .S(N3872), .A(N2050), .B(N3997), .CI(N2813));
ADDFHX1 inst_cellmath__43_0_I1368 (.CO(N3152), .S(N2690), .A(N2958), .B(N3733), .CI(N3872));
ADDFX1 inst_cellmath__43_0_I1369 (.CO(N4066), .S(N3618), .A(N2992), .B(N2771), .CI(N3893));
ADDFXL inst_cellmath__43_0_I1370 (.CO(N2884), .S(N2427), .A(N2421), .B(N3621), .CI(N2705));
ADDFX1 inst_cellmath__43_0_I1371 (.CO(N3795), .S(N3341), .A(N2135), .B(N3040), .CI(N3324));
ADDFX1 inst_cellmath__43_0_I1372 (.CO(N2613), .S(N2164), .A(N3941), .B(N3668), .CI(N2746));
ADDFX1 inst_cellmath__43_0_I1373 (.CO(N3538), .S(N3078), .A(N3373), .B(N2469), .CI(N2182));
ADDFX1 inst_cellmath__43_0_I1374 (.CO(N2347), .S(N3987), .A(N3991), .B(N3091), .CI(N2795));
ADDFXL inst_cellmath__43_0_I1375 (.CO(N3263), .S(N2803), .A(N3467), .B(N3709), .CI(N2281));
ADDFX1 inst_cellmath__43_0_I1376 (.CO(N2085), .S(N3723), .A(N2015), .B(N3197), .CI(N2928));
ADDFXL inst_cellmath__43_0_I1377 (.CO(N2995), .S(N2535), .A(N3838), .B(N3618), .CI(N2427));
ADDFXL inst_cellmath__43_0_I1378 (.CO(N3905), .S(N3458), .A(N2164), .B(N3341), .CI(N3078));
ADDFHXL inst_cellmath__43_0_I1379 (.CO(N2724), .S(N2268), .A(N3987), .B(N2657), .CI(N3585));
ADDFXL inst_cellmath__43_0_I1380 (.CO(N3649), .S(N3188), .A(N2803), .B(N2392), .CI(N3723));
ADDFX1 inst_cellmath__43_0_I1381 (.CO(N2462), .S(N4103), .A(N2125), .B(N3307), .CI(N2535));
ADDFHXL inst_cellmath__43_0_I1382 (.CO(N3377), .S(N2915), .A(N3458), .B(N3039), .CI(N2268));
ADDFHXL inst_cellmath__43_0_I1383 (.CO(N2195), .S(N3828), .A(N2763), .B(N3949), .CI(N3188));
ADDFHXL inst_cellmath__43_0_I1384 (.CO(N3109), .S(N2649), .A(N4103), .B(N3689), .CI(N2915));
ADDFHXL inst_cellmath__43_0_I1385 (.CO(N4020), .S(N3574), .A(N3828), .B(N2504), .CI(N3422));
ADDFHX1 inst_cellmath__43_0_I1386 (.CO(N2834), .S(N2381), .A(N2649), .B(N2233), .CI(N3574));
ADDFX1 inst_cellmath__43_0_I1387 (.CO(N3753), .S(N3297), .A(N2712), .B(N3697), .CI(N3631));
ADDFX1 inst_cellmath__43_0_I1388 (.CO(N2572), .S(N2116), .A(N3335), .B(N2430), .CI(N2147));
ADDFX1 inst_cellmath__43_0_I1389 (.CO(N3492), .S(N3030), .A(N2755), .B(N3047), .CI(N3947));
ADDFXL inst_cellmath__43_0_I1390 (.CO(N2303), .S(N3942), .A(N2475), .B(N3676), .CI(N3383));
ADDFXL inst_cellmath__43_0_I1391 (.CO(N3222), .S(N2756), .A(N3099), .B(N2191), .CI(N4001));
ADDFXL inst_cellmath__43_0_I1392 (.CO(N2040), .S(N3682), .A(N3717), .B(N2805), .CI(N2521));
ADDFX1 inst_cellmath__43_0_I1393 (.CO(N2952), .S(N2495), .A(N4066), .B(N3795), .CI(N2884));
ADDFX1 inst_cellmath__43_0_I1394 (.CO(N3865), .S(N3414), .A(N2613), .B(N3538), .CI(N2347));
ADDFX1 inst_cellmath__43_0_I1395 (.CO(N2681), .S(N2225), .A(N2116), .B(N3030), .CI(N3297));
ADDFXL inst_cellmath__43_0_I1396 (.CO(N3607), .S(N3144), .A(N2756), .B(N3942), .CI(N3682));
ADDFX1 inst_cellmath__43_0_I1397 (.CO(N2419), .S(N4058), .A(N3263), .B(N2085), .CI(N2995));
ADDFX1 inst_cellmath__43_0_I1398 (.CO(N3333), .S(N2874), .A(N2495), .B(N3905), .CI(N3414));
ADDFXL inst_cellmath__43_0_I1399 (.CO(N2153), .S(N3787), .A(N3144), .B(N2724), .CI(N2225));
ADDFXL inst_cellmath__43_0_I1400 (.CO(N3068), .S(N2606), .A(N3649), .B(N2462), .CI(N4058));
ADDFXL inst_cellmath__43_0_I1401 (.CO(N3977), .S(N3528), .A(N3377), .B(N2874), .CI(N3787));
ADDFHXL inst_cellmath__43_0_I1402 (.CO(N2789), .S(N2340), .A(N2606), .B(N2195), .CI(N3109));
ADDFHXL inst_cellmath__43_0_I1403 (.CO(N3716), .S(N3255), .A(N4020), .B(N3528), .CI(N2340));
ADDFXL inst_cellmath__43_0_I1404 (.CO(N2526), .S(N2076), .A(N2512), .B(N2438), .CI(N3344));
ADDFX1 inst_cellmath__43_0_I1405 (.CO(N3450), .S(N2986), .A(N3059), .B(N2159), .CI(N3956));
ADDFX1 inst_cellmath__43_0_I1406 (.CO(N2257), .S(N3897), .A(N3684), .B(N2762), .CI(N2484));
ADDFX1 inst_cellmath__43_0_I1407 (.CO(N3177), .S(N2715), .A(N2200), .B(N3392), .CI(N3108));
ADDFX1 inst_cellmath__43_0_I1408 (.CO(N4092), .S(N3640), .A(N2814), .B(N4007), .CI(N3727));
ADDFX1 inst_cellmath__43_0_I1409 (.CO(N2907), .S(N2452), .A(N3444), .B(N2530), .CI(N3753));
ADDFXL inst_cellmath__43_0_I1410 (.CO(N3818), .S(N3367), .A(N2303), .B(N2572), .CI(N3492));
ADDFX1 inst_cellmath__43_0_I1411 (.CO(N2640), .S(N2187), .A(N2040), .B(N3222), .CI(N2076));
ADDFXL inst_cellmath__43_0_I1412 (.CO(N3563), .S(N3101), .A(N3897), .B(N2986), .CI(N2715));
ADDFX1 inst_cellmath__43_0_I1413 (.CO(N2371), .S(N4012), .A(N3640), .B(N2952), .CI(N3865));
ADDFX1 inst_cellmath__43_0_I1414 (.CO(N3287), .S(N2824), .A(N2452), .B(N3367), .CI(N2681));
ADDFXL inst_cellmath__43_0_I1415 (.CO(N2107), .S(N3744), .A(N3607), .B(N2187), .CI(N3101));
ADDFX1 inst_cellmath__43_0_I1416 (.CO(N3018), .S(N2562), .A(N3333), .B(N2419), .CI(N4012));
ADDFX1 inst_cellmath__43_0_I1417 (.CO(N3933), .S(N3482), .A(N2153), .B(N2824), .CI(N3744));
ADDFXL inst_cellmath__43_0_I1418 (.CO(N2747), .S(N2293), .A(N2562), .B(N3068), .CI(N3977));
ADDFHX1 inst_cellmath__43_0_I1419 (.CO(N3674), .S(N3212), .A(N2789), .B(N3482), .CI(N2293));
ADDFX1 inst_cellmath__43_0_I1420 (.CO(N2485), .S(N2028), .A(N2167), .B(N3431), .CI(N3070));
ADDFX1 inst_cellmath__43_0_I1421 (.CO(N3403), .S(N2942), .A(N3969), .B(N3690), .CI(N2772));
ADDFXL inst_cellmath__43_0_I1422 (.CO(N2216), .S(N3853), .A(N3401), .B(N2493), .CI(N2210));
ADDFX1 inst_cellmath__43_0_I1423 (.CO(N3133), .S(N2672), .A(N4017), .B(N3117), .CI(N2821));
ADDFX1 inst_cellmath__43_0_I1424 (.CO(N4047), .S(N3599), .A(N2540), .B(N3735), .CI(N3452));
ADDFX1 inst_cellmath__43_0_I1425 (.CO(N2865), .S(N2409), .A(N2249), .B(N2526), .CI(N3450));
ADDFX1 inst_cellmath__43_0_I1426 (.CO(N3779), .S(N3322), .A(N3177), .B(N2257), .CI(N4092));
ADDFXL inst_cellmath__43_0_I1427 (.CO(N2598), .S(N2141), .A(N2028), .B(N3853), .CI(N2942));
ADDFXL inst_cellmath__43_0_I1428 (.CO(N3518), .S(N3057), .A(N3599), .B(N2672), .CI(N2907));
ADDFX1 inst_cellmath__43_0_I1429 (.CO(N2331), .S(N3967), .A(N2640), .B(N3818), .CI(N2409));
ADDFXL inst_cellmath__43_0_I1430 (.CO(N3245), .S(N2780), .A(N3322), .B(N3563), .CI(N2141));
ADDFX1 inst_cellmath__43_0_I1431 (.CO(N2067), .S(N3707), .A(N2371), .B(N3057), .CI(N3287));
ADDFX1 inst_cellmath__43_0_I1432 (.CO(N2975), .S(N2516), .A(N2107), .B(N3967), .CI(N2780));
ADDFHXL inst_cellmath__43_0_I1433 (.CO(N3889), .S(N3439), .A(N3018), .B(N3707), .CI(N3933));
ADDFHXL inst_cellmath__43_0_I1434 (.CO(N2706), .S(N2248), .A(N2747), .B(N2516), .CI(N3439));
ADDFX1 inst_cellmath__43_0_I1435 (.CO(N3635), .S(N3168), .A(N3981), .B(N2239), .CI(N2785));
ADDFX1 inst_cellmath__43_0_I1436 (.CO(N2444), .S(N4080), .A(N3413), .B(N3698), .CI(N2503));
ADDFXL inst_cellmath__43_0_I1437 (.CO(N3356), .S(N2899), .A(N3123), .B(N2218), .CI(N4024));
ADDFX1 inst_cellmath__43_0_I1438 (.CO(N2178), .S(N3810), .A(N3743), .B(N2829), .CI(N2550));
ADDFX1 inst_cellmath__43_0_I1439 (.CO(N3092), .S(N2628), .A(N2259), .B(N3459), .CI(N3172));
ADDFX1 inst_cellmath__43_0_I1440 (.CO(N4002), .S(N3554), .A(N3403), .B(N2485), .CI(N2216));
ADDFX1 inst_cellmath__43_0_I1441 (.CO(N2818), .S(N2361), .A(N4047), .B(N3133), .CI(N3168));
ADDFX1 inst_cellmath__43_0_I1442 (.CO(N3736), .S(N3277), .A(N2899), .B(N4080), .CI(N3810));
ADDFX1 inst_cellmath__43_0_I1443 (.CO(N2552), .S(N2096), .A(N2865), .B(N2628), .CI(N3779));
ADDFXL inst_cellmath__43_0_I1444 (.CO(N3470), .S(N3008), .A(N3554), .B(N2598), .CI(N3518));
ADDFX1 inst_cellmath__43_0_I1445 (.CO(N2285), .S(N3923), .A(N3277), .B(N2361), .CI(N2331));
ADDFXL inst_cellmath__43_0_I1446 (.CO(N3204), .S(N2737), .A(N2096), .B(N3245), .CI(N3008));
ADDFX1 inst_cellmath__43_0_I1447 (.CO(N2020), .S(N3666), .A(N3923), .B(N2067), .CI(N2975));
ADDFHXL inst_cellmath__43_0_I1448 (.CO(N2933), .S(N2476), .A(N3889), .B(N2737), .CI(N3666));
ADDFX1 inst_cellmath__43_0_I1449 (.CO(N3845), .S(N3393), .A(N3710), .B(N3162), .CI(N2509));
ADDFXL inst_cellmath__43_0_I1450 (.CO(N2662), .S(N2208), .A(N2227), .B(N3423), .CI(N3131));
ADDFX1 inst_cellmath__43_0_I1451 (.CO(N3590), .S(N3124), .A(N2842), .B(N4033), .CI(N3751));
ADDFX1 inst_cellmath__43_0_I1452 (.CO(N2399), .S(N4034), .A(N3468), .B(N2556), .CI(N2273));
ADDFX1 inst_cellmath__43_0_I1453 (.CO(N3312), .S(N2851), .A(N4084), .B(N3183), .CI(N3635));
ADDFX1 inst_cellmath__43_0_I1454 (.CO(N2130), .S(N3768), .A(N3356), .B(N2444), .CI(N2178));
ADDFX1 inst_cellmath__43_0_I1455 (.CO(N3045), .S(N2587), .A(N3393), .B(N3092), .CI(N2208));
ADDFX1 inst_cellmath__43_0_I1456 (.CO(N3954), .S(N3506), .A(N4034), .B(N3124), .CI(N4002));
ADDFX1 inst_cellmath__43_0_I1457 (.CO(N2767), .S(N2321), .A(N2851), .B(N2818), .CI(N3736));
ADDFX1 inst_cellmath__43_0_I1458 (.CO(N3696), .S(N3234), .A(N2587), .B(N3768), .CI(N2552));
ADDFHXL inst_cellmath__43_0_I1459 (.CO(N2507), .S(N2056), .A(N3470), .B(N3506), .CI(N2321));
ADDFHXL inst_cellmath__43_0_I1460 (.CO(N3428), .S(N2964), .A(N3234), .B(N2285), .CI(N3204));
ADDFX1 inst_cellmath__43_0_I1461 (.CO(N2238), .S(N3879), .A(N2020), .B(N2056), .CI(N2964));
ADDFX1 inst_cellmath__43_0_I1462 (.CO(N3158), .S(N2695), .A(N3432), .B(N4075), .CI(N2234));
ADDFX1 inst_cellmath__43_0_I1463 (.CO(N4070), .S(N3626), .A(N4045), .B(N3142), .CI(N2853));
ADDFX1 inst_cellmath__43_0_I1464 (.CO(N2889), .S(N2433), .A(N2567), .B(N3758), .CI(N3475));
ADDFX1 inst_cellmath__43_0_I1465 (.CO(N3801), .S(N3349), .A(N3192), .B(N2284), .CI(N4094));
ADDFX1 inst_cellmath__43_0_I1466 (.CO(N2619), .S(N2169), .A(N3845), .B(N2901), .CI(N2662));
ADDFX1 inst_cellmath__43_0_I1467 (.CO(N3545), .S(N3083), .A(N2399), .B(N3590), .CI(N2695));
ADDFX1 inst_cellmath__43_0_I1468 (.CO(N2353), .S(N3993), .A(N2433), .B(N3626), .CI(N3349));
ADDFXL inst_cellmath__43_0_I1469 (.CO(N3269), .S(N2809), .A(N2130), .B(N3312), .CI(N3045));
ADDFX1 inst_cellmath__43_0_I1470 (.CO(N2089), .S(N3728), .A(N3083), .B(N2169), .CI(N3954));
ADDFX1 inst_cellmath__43_0_I1471 (.CO(N3001), .S(N2543), .A(N2767), .B(N3993), .CI(N2809));
ADDFHXL inst_cellmath__43_0_I1472 (.CO(N3911), .S(N3462), .A(N3728), .B(N3696), .CI(N2507));
ADDFHXL inst_cellmath__43_0_I1473 (.CO(N2730), .S(N2275), .A(N3428), .B(N2543), .CI(N3462));
ADDFX1 inst_cellmath__43_0_I1474 (.CO(N3656), .S(N3195), .A(N3150), .B(N2890), .CI(N4056));
ADDFX1 inst_cellmath__43_0_I1475 (.CO(N2467), .S(N2012), .A(N3766), .B(N2867), .CI(N2575));
ADDFX1 inst_cellmath__43_0_I1476 (.CO(N3384), .S(N2924), .A(N2291), .B(N3487), .CI(N3201));
ADDFX1 inst_cellmath__43_0_I1477 (.CO(N2201), .S(N3835), .A(N2909), .B(N4104), .CI(N3814));
ADDFX1 inst_cellmath__43_0_I1478 (.CO(N3115), .S(N2654), .A(N4070), .B(N3158), .CI(N2889));
ADDFX1 inst_cellmath__43_0_I1479 (.CO(N4025), .S(N3581), .A(N3195), .B(N3801), .CI(N2012));
ADDFX1 inst_cellmath__43_0_I1480 (.CO(N2840), .S(N2388), .A(N3835), .B(N2924), .CI(N2619));
ADDFX1 inst_cellmath__43_0_I1481 (.CO(N3759), .S(N3302), .A(N2353), .B(N3545), .CI(N2654));
ADDFX1 inst_cellmath__43_0_I1482 (.CO(N2576), .S(N2121), .A(N2388), .B(N3581), .CI(N3269));
ADDFXL inst_cellmath__43_0_I1483 (.CO(N3497), .S(N3038), .A(N3302), .B(N2089), .CI(N3001));
ADDFHX1 inst_cellmath__43_0_I1484 (.CO(N2312), .S(N3945), .A(N3911), .B(N2121), .CI(N3038));
ADDFX1 inst_cellmath__43_0_I1485 (.CO(N3227), .S(N2760), .A(N2876), .B(N3805), .CI(N3777));
ADDFX1 inst_cellmath__43_0_I1486 (.CO(N2045), .S(N3688), .A(N3499), .B(N2585), .CI(N2301));
ADDFX1 inst_cellmath__43_0_I1487 (.CO(N2957), .S(N2500), .A(N2016), .B(N3208), .CI(N2920));
ADDFX1 inst_cellmath__43_0_I1488 (.CO(N3868), .S(N3419), .A(N2633), .B(N3824), .CI(N3656));
ADDFX1 inst_cellmath__43_0_I1489 (.CO(N2687), .S(N2232), .A(N3384), .B(N2467), .CI(N2201));
ADDFX1 inst_cellmath__43_0_I1490 (.CO(N3615), .S(N3147), .A(N3688), .B(N2760), .CI(N2500));
ADDFX1 inst_cellmath__43_0_I1491 (.CO(N2423), .S(N4064), .A(N3419), .B(N3115), .CI(N4025));
ADDFX1 inst_cellmath__43_0_I1492 (.CO(N3338), .S(N2881), .A(N2840), .B(N2232), .CI(N3147));
ADDFX1 inst_cellmath__43_0_I1493 (.CO(N2161), .S(N3792), .A(N4064), .B(N3759), .CI(N2576));
ADDFX1 inst_cellmath__43_0_I1494 (.CO(N3073), .S(N2610), .A(N3497), .B(N2881), .CI(N3792));
ADDFX1 inst_cellmath__43_0_I1495 (.CO(N3984), .S(N3536), .A(N2597), .B(N2623), .CI(N3508));
ADDFX1 inst_cellmath__43_0_I1496 (.CO(N2798), .S(N2345), .A(N3216), .B(N2311), .CI(N2024));
ADDFX1 inst_cellmath__43_0_I1497 (.CO(N3719), .S(N3260), .A(N3832), .B(N2930), .CI(N2642));
ADDFX1 inst_cellmath__43_0_I1498 (.CO(N2531), .S(N2082), .A(N3227), .B(N3556), .CI(N2045));
ADDFX1 inst_cellmath__43_0_I1499 (.CO(N3454), .S(N2993), .A(N3536), .B(N2957), .CI(N2345));
ADDFX1 inst_cellmath__43_0_I1500 (.CO(N2263), .S(N3902), .A(N3868), .B(N3260), .CI(N2687));
ADDFX1 inst_cellmath__43_0_I1501 (.CO(N3185), .S(N2721), .A(N3615), .B(N2082), .CI(N2993));
ADDFX1 inst_cellmath__43_0_I1502 (.CO(N4098), .S(N3646), .A(N3902), .B(N2423), .CI(N3338));
ADDFX1 inst_cellmath__43_0_I1503 (.CO(N2912), .S(N2459), .A(N2161), .B(N2721), .CI(N3646));
ADDFX1 inst_cellmath__43_0_I1504 (.CO(N3826), .S(N3374), .A(N2319), .B(N3546), .CI(N3226));
ADDFX1 inst_cellmath__43_0_I1505 (.CO(N2646), .S(N2193), .A(N2939), .B(N2034), .CI(N3842));
ADDFX1 inst_cellmath__43_0_I1506 (.CO(N3569), .S(N3106), .A(N3565), .B(N2650), .CI(N2366));
ADDFX1 inst_cellmath__43_0_I1507 (.CO(N2379), .S(N4018), .A(N2798), .B(N3984), .CI(N3719));
ADDFX1 inst_cellmath__43_0_I1508 (.CO(N3293), .S(N2831), .A(N2193), .B(N3374), .CI(N3106));
ADDFX1 inst_cellmath__43_0_I1509 (.CO(N2113), .S(N3749), .A(N3454), .B(N2531), .CI(N4018));
ADDFX1 inst_cellmath__43_0_I1510 (.CO(N3027), .S(N2568), .A(N2831), .B(N2263), .CI(N3185));
ADDFX1 inst_cellmath__43_0_I1511 (.CO(N3939), .S(N3489), .A(N4098), .B(N3749), .CI(N2568));
ADDFX1 inst_cellmath__43_0_I1512 (.CO(N2753), .S(N2299), .A(N2047), .B(N2357), .CI(N2950));
ADDFX1 inst_cellmath__43_0_I1513 (.CO(N3680), .S(N3218), .A(N2658), .B(N3849), .CI(N3578));
ADDFX1 inst_cellmath__43_0_I1514 (.CO(N2491), .S(N2036), .A(N3281), .B(N2375), .CI(N3826));
ADDFX1 inst_cellmath__43_0_I1515 (.CO(N3411), .S(N2948), .A(N3569), .B(N2646), .CI(N2299));
ADDFX1 inst_cellmath__43_0_I1516 (.CO(N2222), .S(N3861), .A(N2379), .B(N3218), .CI(N2036));
ADDFX1 inst_cellmath__43_0_I1517 (.CO(N3139), .S(N2677), .A(N2948), .B(N3293), .CI(N2113));
ADDFX1 inst_cellmath__43_0_I1518 (.CO(N4053), .S(N3604), .A(N3027), .B(N3861), .CI(N2677));
ADDFX1 inst_cellmath__43_0_I1519 (.CO(N2873), .S(N2415), .A(N3858), .B(N3274), .CI(N2667));
ADDFX1 inst_cellmath__43_0_I1520 (.CO(N3784), .S(N3330), .A(N2386), .B(N3587), .CI(N3288));
ADDFX1 inst_cellmath__43_0_I1521 (.CO(N2604), .S(N2151), .A(N2753), .B(N2099), .CI(N3680));
ADDFX1 inst_cellmath__43_0_I1522 (.CO(N3527), .S(N3063), .A(N3330), .B(N2415), .CI(N2491));
ADDFX1 inst_cellmath__43_0_I1523 (.CO(N2337), .S(N3974), .A(N2151), .B(N3411), .CI(N2222));
ADDFX1 inst_cellmath__43_0_I1524 (.CO(N3251), .S(N2788), .A(N3139), .B(N3063), .CI(N3974));
ADDFX1 inst_cellmath__43_0_I1525 (.CO(N2075), .S(N3712), .A(N3597), .B(N2090), .CI(N2396));
ADDFX1 inst_cellmath__43_0_I1526 (.CO(N2982), .S(N2522), .A(N2110), .B(N3298), .CI(N3012));
ADDFX1 inst_cellmath__43_0_I1527 (.CO(N3894), .S(N3446), .A(N3784), .B(N2873), .CI(N3712));
ADDFX1 inst_cellmath__43_0_I1528 (.CO(N2713), .S(N2253), .A(N2604), .B(N2522), .CI(N3527));
ADDFX1 inst_cellmath__43_0_I1529 (.CO(N3638), .S(N3173), .A(N2337), .B(N3446), .CI(N2253));
ADDFX1 inst_cellmath__43_0_I1530 (.CO(N2448), .S(N4087), .A(N3308), .B(N3005), .CI(N2119));
ADDFX1 inst_cellmath__43_0_I1531 (.CO(N3365), .S(N2903), .A(N3926), .B(N3023), .CI(N2075));
ADDFX1 inst_cellmath__43_0_I1532 (.CO(N2184), .S(N3815), .A(N4087), .B(N2982), .CI(N3894));
ADDFX1 inst_cellmath__43_0_I1533 (.CO(N3097), .S(N2636), .A(N2713), .B(N2903), .CI(N3815));
ADDFX1 inst_cellmath__43_0_I1534 (.CO(N4009), .S(N3559), .A(N3035), .B(N3915), .CI(N3934));
ADDFX1 inst_cellmath__43_0_I1535 (.CO(N2822), .S(N2369), .A(N2448), .B(N2740), .CI(N3559));
ADDFX1 inst_cellmath__43_0_I1536 (.CO(N3741), .S(N3284), .A(N2369), .B(N3365), .CI(N2184));
ADDFX1 inst_cellmath__43_0_I1537 (.CO(N2558), .S(N2103), .A(N2750), .B(N2731), .CI(N3670));
ADDFX1 inst_cellmath__43_0_I1538 (.CO(N3477), .S(N3015), .A(N2103), .B(N4009), .CI(N2822));
ADDFX1 inst_cellmath__43_0_I1539 (.CO(N2289), .S(N3930), .A(N2478), .B(N3661), .CI(N2558));
OR4X1 inst_cellmath__43_0_I11236 (.Y(N2744), .A(N3075), .B(N3878), .C(N3347), .D(N3614));
NOR2XL inst_cellmath__43_0_I1541 (.Y(N3209), .A(N3752), .B(N2428));
NAND2XL inst_cellmath__43_0_I1542 (.Y(N3672), .A(N3752), .B(N2428));
AND2XL inst_cellmath__43_0_I1544 (.Y(N2482), .A(N3342), .B(N2162));
NOR2XL inst_cellmath__43_0_I1545 (.Y(N2937), .A(N2614), .B(N2799));
NAND2XL inst_cellmath__43_0_I1546 (.Y(N3399), .A(N2614), .B(N2799));
AND2XL inst_cellmath__43_0_I1548 (.Y(N2214), .A(N3455), .B(N2269));
NOR2XL inst_cellmath__43_0_I1549 (.Y(N2669), .A(N2722), .B(N2647));
NAND2XL inst_cellmath__43_0_I1550 (.Y(N3129), .A(N2722), .B(N2647));
AND2XL inst_cellmath__43_0_I1552 (.Y(N4042), .A(N3110), .B(N3940));
NOR2XL inst_cellmath__43_0_I1553 (.Y(N2406), .A(N2304), .B(N4059));
NAND2XL inst_cellmath__43_0_I1554 (.Y(N2862), .A(N2304), .B(N4059));
NOR2XL inst_cellmath__43_0_I1555 (.Y(N3319), .A(N2417), .B(N2987));
NAND2X1 inst_cellmath__43_0_I1556 (.Y(N3775), .A(N2417), .B(N2987));
NOR2XL inst_cellmath__43_0_I1557 (.Y(N2138), .A(N3447), .B(N2825));
NOR2XL inst_cellmath__43_0_I1559 (.Y(N3054), .A(N3285), .B(N3600));
NAND2XL inst_cellmath__43_0_I1560 (.Y(N3516), .A(N3285), .B(N3600));
NOR2XL inst_cellmath__43_0_I1561 (.Y(N3961), .A(N4048), .B(N3169));
NAND2XL inst_cellmath__43_0_I1562 (.Y(N2329), .A(N4048), .B(N3169));
NOR2XL inst_cellmath__43_0_I1563 (.Y(N2777), .A(N3634), .B(N3667));
NAND2X1 inst_cellmath__43_0_I1566 (.Y(N2063), .A(N2021), .B(N2963));
AOI21XL inst_cellmath__43_0_I1567 (.Y(N3435), .A0(N3672), .A1(N2744), .B0(N3209));
OAI22XL inst_cellmath__43_0_I4122 (.Y(N2893), .A0(N2482), .A1(N3435), .B0(N3342), .B1(N2162));
AOI21XL inst_cellmath__43_0_I1571 (.Y(N2358), .A0(N3399), .A1(N2893), .B0(N2937));
OAI22XL inst_cellmath__43_0_I4123 (.Y(N3663), .A0(N2214), .A1(N2358), .B0(N3455), .B1(N2269));
AOI21XL inst_cellmath__43_0_I1575 (.Y(N2847), .A0(N3129), .A1(N3663), .B0(N2669));
OAI22XL inst_cellmath__43_0_I4124 (.Y(N3876), .A0(N4042), .A1(N2847), .B0(N3110), .B1(N3940));
AOI21XL inst_cellmath__43_0_I1579 (.Y(N3623), .A0(N3775), .A1(N2406), .B0(N3319));
INVXL inst_cellmath__43_0_I1580 (.Y(N3916), .A(N3623));
AOI31X1 inst_cellmath__43_0_I1582 (.Y(N3194), .A0(N3775), .A1(N2862), .A2(N3876), .B0(N3916));
AOI21X1 inst_cellmath__43_0_I1583 (.Y(N2918), .A0(N3516), .A1(N2138), .B0(N3054));
OAI2BB1X1 inst_cellmath__43_0_I4125 (.Y(N3380), .A0N(N3447), .A1N(N2825), .B0(N3516));
OAI21X1 inst_cellmath__43_0_I1585 (.Y(N2496), .A0(N3380), .A1(N3194), .B0(N2918));
AOI21X1 inst_cellmath__43_0_I1588 (.Y(N2988), .A0(N2329), .A1(N2496), .B0(N3961));
AOI2BB2X1 inst_cellmath__43_0_I4127 (.Y(N2717), .A0N(N2021), .A1N(N2963), .B0(N2063), .B1(N2777));
OAI2BB1X1 inst_cellmath__43_0_I4128 (.Y(N3181), .A0N(N3634), .A1N(N3667), .B0(N2063));
OAI21X1 inst_cellmath__43_0_I1594 (.Y(N2665), .A0(N3181), .A1(N2988), .B0(N2717));
NOR2XL inst_cellmath__43_0_I1622 (.Y(N3592), .A(N3429), .B(N3196));
NAND2XL inst_cellmath__43_0_I1623 (.Y(N4038), .A(N3429), .B(N3196));
NOR2XL inst_cellmath__43_0_I1624 (.Y(N2402), .A(N3657), .B(N2230));
NOR2XL inst_cellmath__43_0_I1626 (.Y(N3315), .A(N2688), .B(N2194));
NAND2XL inst_cellmath__43_0_I1627 (.Y(N3770), .A(N2688), .B(N2194));
NOR2XL inst_cellmath__43_0_I1628 (.Y(N2136), .A(N2644), .B(N3064));
NAND2X1 inst_cellmath__43_0_I1631 (.Y(N3513), .A(N3523), .B(N2745));
NOR2X1 inst_cellmath__43_0_I1632 (.Y(N3957), .A(N3207), .B(N3354));
NAND2X1 inst_cellmath__43_0_I1633 (.Y(N2324), .A(N3207), .B(N3354));
NOR2XL inst_cellmath__43_0_I1634 (.Y(N2775), .A(N3807), .B(N2764));
NAND2X2 inst_cellmath__43_0_I1635 (.Y(N3237), .A(N3807), .B(N2764));
NOR2X2 inst_cellmath__43_0_I1636 (.Y(N3700), .A(N3233), .B(N4022));
NAND2XL inst_cellmath__43_0_I1637 (.Y(N2061), .A(N3233), .B(N4022));
NOR2X2 inst_cellmath__43_0_I1638 (.Y(N2510), .A(N2385), .B(N3182));
NAND2X4 inst_cellmath__43_0_I1639 (.Y(N2967), .A(N2385), .B(N3182));
NOR2X2 inst_cellmath__43_0_I1640 (.Y(N3433), .A(N3643), .B(N2333));
NAND2X2 inst_cellmath__43_0_I1641 (.Y(N3882), .A(N3643), .B(N2333));
NOR2X2 inst_cellmath__43_0_I1642 (.Y(N2240), .A(N3048), .B(N2783));
NOR2X2 inst_cellmath__43_0_I1644 (.Y(N3160), .A(N3125), .B(N2092));
NAND2X2 inst_cellmath__43_0_I1645 (.Y(N3628), .A(N3125), .B(N2092));
NOR2X1 inst_cellmath__43_0_I1646 (.Y(N4076), .A(N2546), .B(N2690));
NAND2X4 inst_cellmath__43_0_I1647 (.Y(N2436), .A(N2546), .B(N2690));
NOR2X2 inst_cellmath__43_0_I1648 (.Y(N2891), .A(N3152), .B(N2381));
NAND2X4 inst_cellmath__43_0_I1649 (.Y(N3353), .A(N3152), .B(N2381));
NOR2X1 inst_cellmath__43_0_I1650 (.Y(N3803), .A(N2834), .B(N3255));
NAND2X4 inst_cellmath__43_0_I1651 (.Y(N2172), .A(N2834), .B(N3255));
NOR2X2 inst_cellmath__43_0_I1652 (.Y(N2626), .A(N3716), .B(N3212));
NAND2X1 inst_cellmath__43_0_I1653 (.Y(N3087), .A(N3716), .B(N3212));
NOR2X1 inst_cellmath__43_0_I1654 (.Y(N3548), .A(N3674), .B(N2248));
NAND2X4 inst_cellmath__43_0_I1655 (.Y(N3999), .A(N3674), .B(N2248));
NOR2X1 inst_cellmath__43_0_I1656 (.Y(N2355), .A(N2706), .B(N2476));
NAND2X2 inst_cellmath__43_0_I1657 (.Y(N2812), .A(N2706), .B(N2476));
NOR2XL inst_cellmath__43_0_I1658 (.Y(N3275), .A(N2933), .B(N3879));
NAND2X2 inst_cellmath__43_0_I1659 (.Y(N3732), .A(N2933), .B(N3879));
NOR2X2 inst_cellmath__43_0_I1660 (.Y(N2091), .A(N2238), .B(N2275));
NAND2X2 inst_cellmath__43_0_I1661 (.Y(N2548), .A(N2238), .B(N2275));
NOR2X1 inst_cellmath__43_0_I1662 (.Y(N3003), .A(N2730), .B(N3945));
NAND2X4 inst_cellmath__43_0_I1663 (.Y(N3466), .A(N2730), .B(N3945));
NOR2XL inst_cellmath__43_0_I1664 (.Y(N3917), .A(N2312), .B(N2610));
NAND2X1 inst_cellmath__43_0_I1665 (.Y(N2280), .A(N2312), .B(N2610));
NOR2XL inst_cellmath__43_0_I1666 (.Y(N2732), .A(N3073), .B(N2459));
NAND2X1 inst_cellmath__43_0_I1667 (.Y(N3199), .A(N3073), .B(N2459));
NOR2XL inst_cellmath__43_0_I1668 (.Y(N3659), .A(N2912), .B(N3489));
NAND2XL inst_cellmath__43_0_I1669 (.Y(N2014), .A(N2912), .B(N3489));
NOR2XL inst_cellmath__43_0_I1670 (.Y(N2471), .A(N3939), .B(N3604));
NAND2XL inst_cellmath__43_0_I1671 (.Y(N2927), .A(N3939), .B(N3604));
NOR2XL inst_cellmath__43_0_I1672 (.Y(N3386), .A(N4053), .B(N2788));
NAND2XL inst_cellmath__43_0_I1673 (.Y(N3840), .A(N4053), .B(N2788));
NOR2XL inst_cellmath__43_0_I1674 (.Y(N2203), .A(N3251), .B(N3173));
NAND2XL inst_cellmath__43_0_I1675 (.Y(N2656), .A(N3251), .B(N3173));
NOR2XL inst_cellmath__43_0_I1676 (.Y(N3119), .A(N3638), .B(N2636));
NAND2XL inst_cellmath__43_0_I1677 (.Y(N3584), .A(N3638), .B(N2636));
NOR2XL inst_cellmath__43_0_I1678 (.Y(N4028), .A(N3284), .B(N3097));
NAND2XL inst_cellmath__43_0_I1679 (.Y(N2394), .A(N3284), .B(N3097));
NOR2XL inst_cellmath__43_0_I1680 (.Y(N2844), .A(N3015), .B(N3741));
NAND2XL inst_cellmath__43_0_I1681 (.Y(N3306), .A(N3015), .B(N3741));
NOR2XL inst_cellmath__43_0_I1682 (.Y(N3762), .A(N3930), .B(N3477));
NAND2XL inst_cellmath__43_0_I1683 (.Y(N2124), .A(N3930), .B(N3477));
AOI21X1 inst_cellmath__43_0_I1685 (.Y(N3948), .A0(N4038), .A1(N2665), .B0(N3592));
AOI21XL inst_cellmath__43_0_I1686 (.Y(N3691), .A0(N3770), .A1(N2402), .B0(N3315));
OAI2BB1X1 inst_cellmath__43_0_I4132 (.Y(N2049), .A0N(N3657), .A1N(N2230), .B0(N3770));
OAI21X1 inst_cellmath__43_0_I1688 (.Y(N3151), .A0(N2049), .A1(N3948), .B0(N3691));
AOI2BB2X1 inst_cellmath__43_0_I4133 (.Y(N2883), .A0N(N3523), .A1N(N2745), .B0(N3513), .B1(N2136));
OAI2BB1X1 inst_cellmath__43_0_I4134 (.Y(N3343), .A0N(N2644), .A1N(N3064), .B0(N3513));
AOI21X1 inst_cellmath__43_0_I1692 (.Y(N2615), .A0(N3237), .A1(N3957), .B0(N2775));
NAND2X2 inst_cellmath__43_0_I1693 (.Y(N3077), .A(N3237), .B(N2324));
OAI21X2 inst_cellmath__43_0_I1694 (.Y(N2084), .A0(N3077), .A1(N2883), .B0(N2615));
NOR2X2 inst_cellmath__43_0_I1695 (.Y(N2538), .A(N3077), .B(N3343));
AOI21X4 inst_cellmath__43_0_I1696 (.Y(N3907), .A0(N3700), .A1(N2967), .B0(N2510));
NAND2X2 inst_cellmath__43_0_I1697 (.Y(N2267), .A(N2967), .B(N2061));
INVXL inst_cellmath__43_0_I1698 (.Y(N2725), .A(N3882));
AOI21X4 inst_cellmath__43_0_I1699 (.Y(N3648), .A0(N3433), .A1(N2701), .B0(N2240));
NAND2X4 inst_cellmath__43_0_I1700 (.Y(N4102), .A(N2701), .B(N3882));
OAI21X4 inst_cellmath__43_0_I1701 (.Y(N3111), .A0(N4102), .A1(N3907), .B0(N3648));
NOR2X2 inst_cellmath__43_0_I1704 (.Y(N3573), .A(N4102), .B(N2267));
AOI21X4 inst_cellmath__43_0_I1705 (.Y(N2833), .A0(N3160), .A1(N2436), .B0(N4076));
NAND2X4 inst_cellmath__43_0_I1706 (.Y(N3296), .A(N3628), .B(N2436));
INVXL inst_cellmath__43_0_I1707 (.Y(N2836), .A(N3353));
AOI21X4 inst_cellmath__43_0_I1708 (.Y(N2571), .A0(N2891), .A1(N2172), .B0(N3803));
NAND2X6 inst_cellmath__43_0_I1709 (.Y(N3033), .A(N2172), .B(N3353));
OAI21X4 inst_cellmath__43_0_I1710 (.Y(N2039), .A0(N3033), .A1(N2833), .B0(N2571));
NOR2X6 inst_cellmath__43_0_I1711 (.Y(N2494), .A(N3296), .B(N3033));
AOI21X4 inst_cellmath__43_0_I1712 (.Y(N3864), .A0(N3999), .A1(N2626), .B0(N3548));
NAND2X4 inst_cellmath__43_0_I1713 (.Y(N2228), .A(N3999), .B(N3087));
INVXL inst_cellmath__43_0_I1714 (.Y(N3223), .A(N2812));
AOI21X2 inst_cellmath__43_0_I1715 (.Y(N3609), .A0(N3732), .A1(N2355), .B0(N3275));
NAND2X4 inst_cellmath__43_0_I1716 (.Y(N4057), .A(N3732), .B(N2812));
OAI21X4 inst_cellmath__43_0_I1717 (.Y(N3067), .A0(N4057), .A1(N3864), .B0(N3609));
NOR2X4 inst_cellmath__43_0_I1718 (.Y(N3531), .A(N4057), .B(N2228));
AOI21X4 inst_cellmath__43_0_I1719 (.Y(N2793), .A0(N3466), .A1(N2091), .B0(N3003));
NAND2X2 inst_cellmath__43_0_I1720 (.Y(N3254), .A(N3466), .B(N2548));
INVXL inst_cellmath__43_0_I1721 (.Y(N2683), .A(N2280));
AOI21X1 inst_cellmath__43_0_I1722 (.Y(N2525), .A0(N3917), .A1(N3199), .B0(N2732));
NAND2X2 inst_cellmath__43_0_I1723 (.Y(N2985), .A(N3199), .B(N2280));
OAI21X4 inst_cellmath__43_0_I1724 (.Y(N4091), .A0(N2985), .A1(N2793), .B0(N2525));
NOR2X1 inst_cellmath__43_0_I1725 (.Y(N2454), .A(N2985), .B(N3254));
AOI21XL inst_cellmath__43_0_I1726 (.Y(N3822), .A0(N2927), .A1(N3659), .B0(N2471));
NAND2XL inst_cellmath__43_0_I1727 (.Y(N2186), .A(N2927), .B(N2014));
INVXL inst_cellmath__43_0_I1728 (.Y(N3788), .A(N3386));
INVXL inst_cellmath__43_0_I1729 (.Y(N2156), .A(N3840));
AOI21XL inst_cellmath__43_0_I1730 (.Y(N3562), .A0(N2656), .A1(N3386), .B0(N2203));
NAND2XL inst_cellmath__43_0_I1731 (.Y(N4011), .A(N2656), .B(N3840));
INVXL inst_cellmath__43_0_I1732 (.Y(N3530), .A(N3822));
INVXL inst_cellmath__43_0_I1733 (.Y(N3979), .A(N2186));
OAI21XL inst_cellmath__43_0_I1734 (.Y(N2106), .A0(N2156), .A1(N3822), .B0(N3788));
NOR2XL inst_cellmath__43_0_I1735 (.Y(N2561), .A(N2156), .B(N2186));
OAI21XL inst_cellmath__43_0_I1736 (.Y(N3021), .A0(N4011), .A1(N3822), .B0(N3562));
NOR2XL inst_cellmath__43_0_I1737 (.Y(N3481), .A(N4011), .B(N2186));
AOI21XL inst_cellmath__43_0_I1738 (.Y(N3402), .A0(N2014), .A1(N4091), .B0(N3659));
AOI21XL inst_cellmath__43_0_I1739 (.Y(N2219), .A0(N3979), .A1(N4091), .B0(N3530));
AOI21XL inst_cellmath__43_0_I1740 (.Y(N3132), .A0(N2561), .A1(N4091), .B0(N2106));
AOI21X2 inst_cellmath__43_0_I1741 (.Y(N4046), .A0(N3481), .A1(N4091), .B0(N3021));
AOI21XL inst_cellmath__43_0_I1742 (.Y(N3778), .A0(N2394), .A1(N3119), .B0(N4028));
NAND2XL inst_cellmath__43_0_I1743 (.Y(N2144), .A(N2394), .B(N3584));
INVXL inst_cellmath__43_0_I1744 (.Y(N3180), .A(N3306));
AOI21XL inst_cellmath__43_0_I1745 (.Y(N3520), .A0(N2124), .A1(N2844), .B0(N3762));
NAND2XL inst_cellmath__43_0_I1746 (.Y(N3966), .A(N2124), .B(N3306));
INVX1 inst_cellmath__43_0_I1751 (.Y(N2944), .A(N4046));
CLKAND2X2 inst_cellmath__43_0_I1752 (.Y(N3405), .A(N3481), .B(N2454));
INVXL inst_cellmath__43_0_I1753 (.Y(N2143), .A(N3151));
AOI21X1 inst_cellmath__43_0_I1755 (.Y(N3767), .A0(N3573), .A1(N2084), .B0(N3111));
NAND2X1 inst_cellmath__43_0_I1756 (.Y(N2132), .A(N3573), .B(N2538));
AOI21X1 inst_cellmath__43_0_I1759 (.Y(N3510), .A0(N3531), .A1(N2039), .B0(N3067));
NAND2X2 inst_cellmath__43_0_I1760 (.Y(N3953), .A(N3531), .B(N2494));
INVXL inst_cellmath__43_0_I1763 (.Y(N2332), .A(N2143));
OAI21X2 inst_cellmath__43_0_I1765 (.Y(N2697), .A0(N3953), .A1(N3767), .B0(N3510));
NOR2X2 inst_cellmath__43_0_I1766 (.Y(N3157), .A(N3953), .B(N2132));
AOI21X2 inst_cellmath__43_0_I11204 (.Y(N2854), .A0(N2538), .A1(N3151), .B0(N2084));
INVX2 inst_cellmath__43_0_I11210 (.Y(N2782), .A(N2854));
INVXL inst_cellmath__43_0_I1770 (.Y(N3708), .A(N2782));
OA21X1 inst_cellmath__43_0_I1771 (.Y(N2069), .A0(N2132), .A1(N2143), .B0(N3767));
NAND2X4 inst_cellmath__43_0_I11206 (.Y(N3044), .A(N2494), .B(N3573));
AOI21X4 inst_cellmath__43_0_I11205 (.Y(N2586), .A0(N2494), .A1(N3111), .B0(N2039));
OA21X1 inst_cellmath__43_0_I1772 (.Y(N2518), .A0(N3044), .A1(N2854), .B0(N2586));
AOI21X4 inst_cellmath__43_0_I1773 (.Y(N3995), .A0(N3157), .A1(N2332), .B0(N2697));
AOI21X4 inst_cellmath__43_0_I11207 (.Y(N18901), .A0(N3405), .A1(N3067), .B0(N2944));
NAND2X4 inst_cellmath__43_0_I11208 (.Y(N18886), .A(N3531), .B(N3405));
NOR2X8 inst_cellmath__43_0_I11209 (.Y(N18904), .A(N18886), .B(N3044));
OAI21X4 inst_cellmath__43_0_I11211 (.Y(N18898), .A0(N18886), .A1(N2586), .B0(N18901));
AOI21X2 inst_cellmath__43_0_I11212 (.Y(N3441), .A0(N18904), .A1(N2782), .B0(N18898));
AOI21X4 inst_cellmath__43_0_I11213 (.Y(N2808), .A0(N2782), .A1(N18904), .B0(N18898));
NOR2XL inst_cellmath__43_0_I1781 (.Y(N2277), .A(N2725), .B(N3907));
NOR2XL inst_cellmath__43_0_I1782 (.Y(N3555), .A(N2277), .B(N3433));
NOR2XL inst_cellmath__43_0_I1783 (.Y(N3385), .A(N2836), .B(N2833));
NOR2XL inst_cellmath__43_0_I1784 (.Y(N2098), .A(N3385), .B(N2891));
NOR2X1 inst_cellmath__43_0_I1785 (.Y(N2391), .A(N3223), .B(N3864));
NOR2XL inst_cellmath__43_0_I1786 (.Y(N2739), .A(N2391), .B(N2355));
NOR2XL inst_cellmath__43_0_I1787 (.Y(N3500), .A(N2683), .B(N2793));
NOR2XL inst_cellmath__43_0_I1788 (.Y(N3395), .A(N3500), .B(N3917));
INVXL inst_cellmath__43_0_I1789 (.Y(N2211), .A(N4091));
NOR2XL inst_cellmath__43_0_I1790 (.Y(N2502), .A(N3180), .B(N3778));
NOR2XL inst_cellmath__43_0_I1791 (.Y(N3509), .A(N2502), .B(N2844));
OAI21XL inst_cellmath__43_0_I11161 (.Y(N2974), .A0(N3966), .A1(N3778), .B0(N3520));
INVXL inst_cellmath__43_0_I1792 (.Y(N2322), .A(N2974));
NAND2BXL inst_cellmath__43_0_I1801 (.Y(N2252), .AN(N2510), .B(N2967));
NAND2BXL inst_cellmath__43_0_I1802 (.Y(N2858), .AN(N3433), .B(N3882));
NAND2BXL inst_cellmath__43_0_I1803 (.Y(N3699), .AN(N2240), .B(N2701));
NAND2BXL inst_cellmath__43_0_I1804 (.Y(N2183), .AN(N3160), .B(N3628));
NAND2BXL inst_cellmath__43_0_I1805 (.Y(N3558), .AN(N4076), .B(N2436));
NAND2BXL inst_cellmath__43_0_I1806 (.Y(N3547), .AN(N2891), .B(N3353));
NAND2BXL inst_cellmath__43_0_I1807 (.Y(N2282), .AN(N3803), .B(N2172));
NAND2BXL inst_cellmath__43_0_I1808 (.Y(N3476), .AN(N2626), .B(N3087));
NAND2BXL inst_cellmath__43_0_I1809 (.Y(N2743), .AN(N3548), .B(N3999));
NAND2BXL inst_cellmath__43_0_I1810 (.Y(N2126), .AN(N2355), .B(N2812));
NAND2BXL inst_cellmath__43_0_I1811 (.Y(N2960), .AN(N3275), .B(N3732));
NAND2BXL inst_cellmath__43_0_I1812 (.Y(N2668), .AN(N2091), .B(N2548));
NAND2BXL inst_cellmath__43_0_I1813 (.Y(N4041), .AN(N3003), .B(N3466));
NAND2BXL inst_cellmath__43_0_I1814 (.Y(N2802), .AN(N3917), .B(N2280));
NAND2BXL inst_cellmath__43_0_I1815 (.Y(N3651), .AN(N2732), .B(N3199));
NAND2BXL inst_cellmath__43_0_I1816 (.Y(N2384), .AN(N3659), .B(N2014));
NAND2BXL inst_cellmath__43_0_I1817 (.Y(N3221), .AN(N2471), .B(N2927));
NAND2BXL inst_cellmath__43_0_I1818 (.Y(N4060), .AN(N3386), .B(N3840));
NAND2BXL inst_cellmath__43_0_I1819 (.Y(N2792), .AN(N2203), .B(N2656));
NAND2BXL inst_cellmath__43_0_I1820 (.Y(N3164), .AN(N3119), .B(N3584));
NAND2BXL inst_cellmath__43_0_I1821 (.Y(N2443), .AN(N4028), .B(N2394));
NAND2BXL inst_cellmath__43_0_I1822 (.Y(N2639), .AN(N2844), .B(N3306));
NAND2BXL inst_cellmath__43_0_I1823 (.Y(N3484), .AN(N3762), .B(N2124));
XNOR2X1 inst_cellmath__43_0_I1830 (.Y(inst_cellmath__43[26]), .A(N2183), .B(N2069));
XNOR2X1 inst_cellmath__43_0_I1831 (.Y(inst_cellmath__43[30]), .A(N2518), .B(N3476));
INVX2 inst_cellmath__43_0_I1832 (.Y(N3149), .A(N3995));
MXI2X1 inst_cellmath__43_0_I1833 (.Y(inst_cellmath__43[34]), .A(N3995), .B(N3149), .S0(N2668));
XNOR2X1 inst_cellmath__43_0_I11242 (.Y(inst_cellmath__43[42]), .A(N3441), .B(N3164));
XNOR2X1 inst_cellmath__43_0_I1846 (.Y(N4031), .A(N2252), .B(N2061));
XNOR2X1 inst_cellmath__43_0_I1847 (.Y(N3588), .A(N3700), .B(N2252));
MXI2XL inst_cellmath__43_0_I1848 (.Y(inst_cellmath__43[23]), .A(N4031), .B(N3588), .S0(N3708));
XOR2XL inst_cellmath__43_0_I1849 (.Y(N2850), .A(N3907), .B(N2858));
NAND2XL inst_cellmath__43_0_I1850 (.Y(N4037), .A(N2267), .B(N3907));
XNOR2X1 inst_cellmath__43_0_I1851 (.Y(N3309), .A(N2858), .B(N4037));
MXI2XL inst_cellmath__43_0_I1852 (.Y(inst_cellmath__43[24]), .A(N3309), .B(N2850), .S0(N3708));
XOR2XL inst_cellmath__43_0_I1853 (.Y(N2128), .A(N3699), .B(N3555));
OAI21XL inst_cellmath__43_0_I1854 (.Y(N2774), .A0(N2725), .A1(N2267), .B0(N3555));
INVXL xnor2_A_I11273 (.Y(N18917), .A(N3699));
MXI2XL xnor2_A_I11274 (.Y(N2583), .A(N3699), .B(N18917), .S0(N2774));
MXI2XL inst_cellmath__43_0_I1856 (.Y(inst_cellmath__43[25]), .A(N2583), .B(N2128), .S0(N3708));
XNOR2X1 inst_cellmath__43_0_I1857 (.Y(N3950), .A(N3628), .B(N3558));
XNOR2X1 inst_cellmath__43_0_I1858 (.Y(N3505), .A(N3160), .B(N3558));
MXI2XL inst_cellmath__43_0_I1859 (.Y(inst_cellmath__43[27]), .A(N3950), .B(N3505), .S0(N2069));
XOR2XL inst_cellmath__43_0_I1860 (.Y(N2765), .A(N2833), .B(N3547));
NAND2XL inst_cellmath__43_0_I1861 (.Y(N2625), .A(N3296), .B(N2833));
XNOR2X1 inst_cellmath__43_0_I1862 (.Y(N3232), .A(N3547), .B(N2625));
MXI2XL inst_cellmath__43_0_I1863 (.Y(inst_cellmath__43[28]), .A(N3232), .B(N2765), .S0(N2069));
XOR2XL inst_cellmath__43_0_I1864 (.Y(N2055), .A(N2282), .B(N2098));
OAI21XL inst_cellmath__43_0_I1865 (.Y(N3465), .A0(N2836), .A1(N3296), .B0(N2098));
INVXL xnor2_A_I11275 (.Y(N18923), .A(N2282));
MXI2XL xnor2_A_I11276 (.Y(N2505), .A(N2282), .B(N18923), .S0(N3465));
MXI2XL inst_cellmath__43_0_I1867 (.Y(inst_cellmath__43[29]), .A(N2505), .B(N2055), .S0(N2069));
XNOR2X1 inst_cellmath__43_0_I1868 (.Y(N3875), .A(N3087), .B(N2743));
XNOR2X1 inst_cellmath__43_0_I1869 (.Y(N3426), .A(N2743), .B(N2626));
MXI2XL inst_cellmath__43_0_I1870 (.Y(inst_cellmath__43[31]), .A(N3875), .B(N3426), .S0(N2518));
XOR2XL inst_cellmath__43_0_I1871 (.Y(N2694), .A(N2126), .B(N3864));
NAND2XL inst_cellmath__43_0_I1872 (.Y(N3305), .A(N2228), .B(N3864));
XNOR2X1 inst_cellmath__43_0_I1873 (.Y(N3154), .A(N2126), .B(N3305));
MXI2XL inst_cellmath__43_0_I1874 (.Y(inst_cellmath__43[32]), .A(N3154), .B(N2694), .S0(N2518));
XOR2XL inst_cellmath__43_0_I1875 (.Y(N4068), .A(N2960), .B(N2739));
OAI21XL inst_cellmath__43_0_I1876 (.Y(N2051), .A0(N3223), .A1(N2228), .B0(N2739));
XNOR2X1 inst_cellmath__43_0_I1877 (.Y(N2431), .A(N2960), .B(N2051));
MXI2XL inst_cellmath__43_0_I1878 (.Y(inst_cellmath__43[33]), .A(N2431), .B(N4068), .S0(N2518));
XNOR2X1 inst_cellmath__43_0_I1879 (.Y(N3797), .A(N4041), .B(N2548));
XNOR2X1 inst_cellmath__43_0_I1880 (.Y(N3348), .A(N4041), .B(N2091));
MXI2XL inst_cellmath__43_0_I1881 (.Y(inst_cellmath__43[35]), .A(N3797), .B(N3348), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1882 (.Y(N2617), .A(N2802), .B(N2793));
NAND2XL inst_cellmath__43_0_I1883 (.Y(N3989), .A(N3254), .B(N2793));
XNOR2X1 inst_cellmath__43_0_I1884 (.Y(N3081), .A(N2802), .B(N3989));
MXI2XL inst_cellmath__43_0_I1885 (.Y(inst_cellmath__43[36]), .A(N3081), .B(N2617), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1886 (.Y(N3992), .A(N3651), .B(N3395));
OAI21XL inst_cellmath__43_0_I1887 (.Y(N2723), .A0(N2683), .A1(N3254), .B0(N3395));
XNOR2X1 inst_cellmath__43_0_I1888 (.Y(N2349), .A(N3651), .B(N2723));
MXI2XL inst_cellmath__43_0_I1889 (.Y(inst_cellmath__43[37]), .A(N2349), .B(N3992), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1890 (.Y(N3267), .A(N2384), .B(N2211));
NAND2BXL inst_cellmath__43_0_I1891 (.Y(N3576), .AN(N2454), .B(N2211));
XNOR2X1 inst_cellmath__43_0_I1892 (.Y(N3725), .A(N2384), .B(N3576));
MXI2XL inst_cellmath__43_0_I1893 (.Y(inst_cellmath__43[38]), .A(N3725), .B(N3267), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1894 (.Y(N2541), .A(N3221), .B(N3402));
OAI2BB1X1 inst_cellmath__43_0_I1895 (.Y(N2305), .A0N(N2014), .A1N(N2454), .B0(N3402));
XNOR2X1 inst_cellmath__43_0_I1896 (.Y(N2997), .A(N3221), .B(N2305));
MXI2XL inst_cellmath__43_0_I1897 (.Y(inst_cellmath__43[39]), .A(N2997), .B(N2541), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1898 (.Y(N3910), .A(N4060), .B(N2219));
OAI2BB1X1 inst_cellmath__43_0_I1899 (.Y(N3143), .A0N(N3979), .A1N(N2454), .B0(N2219));
XNOR2X1 inst_cellmath__43_0_I1900 (.Y(N2270), .A(N4060), .B(N3143));
MXI2XL inst_cellmath__43_0_I1901 (.Y(inst_cellmath__43[40]), .A(N2270), .B(N3910), .S0(N3995));
XOR2XL inst_cellmath__43_0_I1902 (.Y(N3193), .A(N2792), .B(N3132));
OAI2BB1X1 inst_cellmath__43_0_I1903 (.Y(N3980), .A0N(N2561), .A1N(N2454), .B0(N3132));
XNOR2X1 inst_cellmath__43_0_I1904 (.Y(N3654), .A(N2792), .B(N3980));
MXI2XL inst_cellmath__43_0_I1905 (.Y(inst_cellmath__43[41]), .A(N3654), .B(N3193), .S0(N3995));
XNOR2X1 inst_cellmath__43_0_I1906 (.Y(N2922), .A(N2443), .B(N3584));
XNOR2X1 inst_cellmath__43_0_I1907 (.Y(N2466), .A(N2443), .B(N3119));
MXI2XL inst_cellmath__43_0_I1908 (.Y(inst_cellmath__43[43]), .A(N2922), .B(N2466), .S0(N3441));
XOR2XL inst_cellmath__43_0_I1909 (.Y(N3834), .A(N2639), .B(N3778));
NAND2XL inst_cellmath__43_0_I1910 (.Y(N3821), .A(N2144), .B(N3778));
XNOR2X1 inst_cellmath__43_0_I1911 (.Y(N2199), .A(N2639), .B(N3821));
MXI2XL inst_cellmath__43_0_I1912 (.Y(inst_cellmath__43[44]), .A(N2199), .B(N3834), .S0(N3441));
XOR2XL inst_cellmath__43_0_I1913 (.Y(N3114), .A(N3484), .B(N3509));
OAI21XL inst_cellmath__43_0_I1914 (.Y(N2560), .A0(N3180), .A1(N2144), .B0(N3509));
XNOR2X1 inst_cellmath__43_0_I1915 (.Y(N3579), .A(N3484), .B(N2560));
MXI2XL inst_cellmath__43_0_I1916 (.Y(inst_cellmath__43[45]), .A(N3579), .B(N3114), .S0(N3441));
INVXL inst_cellmath__43_0_I11160 (.Y(N2579), .A(N2289));
XNOR2X1 inst_cellmath__43_0_I1917 (.Y(N2387), .A(N2579), .B(N2322));
NOR2XL inst_cellmath__43_0_I11162 (.Y(N3442), .A(N3966), .B(N2144));
NAND2BXL inst_cellmath__43_0_I1918 (.Y(N3406), .AN(N3442), .B(N2322));
XOR2XL inst_cellmath__43_0_I1919 (.Y(N2839), .A(N2579), .B(N3406));
MXI2XL inst_cellmath__43_0_I1920 (.Y(inst_cellmath__43[46]), .A(N2839), .B(N2387), .S0(N3441));
AND2XL inst_cellmath__43_0_I11243 (.Y(N18785), .A(N2579), .B(N2974));
NAND2X2 inst_cellmath__43_0_I11165 (.Y(N18795), .A(N3442), .B(N2579));
NOR2X4 inst_cellmath__43_0_I11170 (.Y(N18799), .A(N18795), .B(N2808));
NOR2X4 inst_cellmath__43_0_I11171 (.Y(inst_cellmath__43[47]), .A(N18785), .B(N18799));
NOR2XL cynw_cm_float_mul_I1922 (.Y(N6156), .A(inst_cellmath__26), .B(inst_cellmath__22));
NOR2XL inst_cellmath__30__14__I1924 (.Y(N6163), .A(inst_cellmath__25), .B(inst_cellmath__21));
NAND2XL inst_cellmath__30__14__I1925 (.Y(N272), .A(N6163), .B(inst_cellmath__24));
OAI2BB1X1 cynw_cm_float_mul_I4143 (.Y(N6169), .A0N(N6156), .A1N(inst_cellmath__23), .B0(N272));
INVXL inst_cellmath__34_0_I1928 (.Y(N6189), .A(a_exp[7]));
INVXL inst_cellmath__34_0_I1929 (.Y(N6263), .A(a_exp[0]));
INVXL inst_cellmath__34_0_I1930 (.Y(N6218), .A(b_exp[0]));
NOR2XL inst_cellmath__34_0_I1931 (.Y(N6176), .A(a_exp[1]), .B(b_exp[1]));
NAND2XL inst_cellmath__34_0_I1932 (.Y(N6254), .A(a_exp[1]), .B(b_exp[1]));
NOR2XL inst_cellmath__34_0_I1933 (.Y(N6184), .A(a_exp[2]), .B(b_exp[2]));
NAND2XL inst_cellmath__34_0_I1934 (.Y(N6204), .A(a_exp[2]), .B(b_exp[2]));
NOR2XL inst_cellmath__34_0_I1935 (.Y(N6227), .A(a_exp[3]), .B(b_exp[3]));
NAND2XL inst_cellmath__34_0_I1936 (.Y(N6240), .A(a_exp[3]), .B(b_exp[3]));
NOR2XL inst_cellmath__34_0_I1937 (.Y(N6259), .A(a_exp[4]), .B(b_exp[4]));
NAND2XL inst_cellmath__34_0_I1938 (.Y(N6193), .A(a_exp[4]), .B(b_exp[4]));
NOR2XL inst_cellmath__34_0_I1939 (.Y(N6213), .A(a_exp[5]), .B(b_exp[5]));
NAND2XL inst_cellmath__34_0_I1940 (.Y(N6232), .A(a_exp[5]), .B(b_exp[5]));
NOR2XL inst_cellmath__34_0_I1941 (.Y(N6249), .A(a_exp[6]), .B(b_exp[6]));
NAND2XL inst_cellmath__34_0_I1942 (.Y(N6180), .A(a_exp[6]), .B(b_exp[6]));
NOR2XL inst_cellmath__34_0_I1943 (.Y(N6201), .A(b_exp[7]), .B(N6189));
NAND2XL inst_cellmath__34_0_I1944 (.Y(N6224), .A(b_exp[7]), .B(N6189));
AND2XL inst_cellmath__34_0_I1945 (.Y(N6210), .A(N6218), .B(N6263));
AND2XL inst_cellmath__34_0_I1946 (.Y(N6237), .A(N6254), .B(N6218));
INVXL inst_cellmath__34_0_I1947 (.Y(N6247), .A(N6184));
OAI2BB1X1 inst_cellmath__34_0_I1948 (.Y(N6256), .A0N(N6204), .A1N(N6176), .B0(N6247));
AND2XL inst_cellmath__34_0_I1949 (.Y(N6186), .A(N6204), .B(N6254));
AO21XL inst_cellmath__34_0_I1950 (.Y(N6206), .A0(N6240), .A1(N6184), .B0(N6227));
AND2XL inst_cellmath__34_0_I1951 (.Y(N6229), .A(N6240), .B(N6204));
AO21XL inst_cellmath__34_0_I1952 (.Y(N6242), .A0(N6193), .A1(N6227), .B0(N6259));
AND2XL inst_cellmath__34_0_I1953 (.Y(N6261), .A(N6193), .B(N6240));
AO21XL inst_cellmath__34_0_I1954 (.Y(N6196), .A0(N6232), .A1(N6259), .B0(N6213));
AND2XL inst_cellmath__34_0_I1955 (.Y(N6215), .A(N6232), .B(N6193));
AO21XL inst_cellmath__34_0_I1956 (.Y(N6233), .A0(N6180), .A1(N6213), .B0(N6249));
AND2XL inst_cellmath__34_0_I1957 (.Y(N6251), .A(N6180), .B(N6232));
AO21XL inst_cellmath__34_0_I1958 (.Y(N6181), .A0(N6224), .A1(N6249), .B0(N6201));
AND2XL inst_cellmath__34_0_I1959 (.Y(N6202), .A(N6224), .B(N6180));
AND2XL inst_cellmath__34_0_I1960 (.Y(N6258), .A(N6189), .B(N6224));
AO21XL inst_cellmath__34_0_I1961 (.Y(N6178), .A0(N6263), .A1(N6237), .B0(N6176));
AO21XL inst_cellmath__34_0_I1962 (.Y(N6222), .A0(N6210), .A1(N6186), .B0(N6256));
AO21XL inst_cellmath__34_0_I1963 (.Y(N6257), .A0(N6176), .A1(N6229), .B0(N6206));
AND2XL inst_cellmath__34_0_I1964 (.Y(N6188), .A(N6229), .B(N6237));
AO21XL inst_cellmath__34_0_I1965 (.Y(N6207), .A0(N6261), .A1(N6256), .B0(N6242));
AND2XL inst_cellmath__34_0_I1966 (.Y(N6230), .A(N6261), .B(N6186));
AO21XL inst_cellmath__34_0_I1967 (.Y(N6244), .A0(N6215), .A1(N6206), .B0(N6196));
AO21XL inst_cellmath__34_0_I1969 (.Y(N6198), .A0(N6251), .A1(N6242), .B0(N6233));
AO21XL inst_cellmath__34_0_I1971 (.Y(N6234), .A0(N6202), .A1(N6196), .B0(N6181));
AND2XL inst_cellmath__34_0_I1972 (.Y(N6253), .A(N6202), .B(N6215));
AO22XL inst_cellmath__34_0_I1973 (.Y(N6183), .A0(N6189), .A1(N6201), .B0(N6258), .B1(N6233));
AND2XL inst_cellmath__34_0_I1974 (.Y(N6203), .A(N6258), .B(N6251));
AO21XL inst_cellmath__34_0_I1975 (.Y(N6175), .A0(N6253), .A1(N6257), .B0(N6234));
AND2XL inst_cellmath__34_0_I1976 (.Y(N6199), .A(N6253), .B(N6188));
AO21XL inst_cellmath__34_0_I1977 (.Y(N6220), .A0(N6203), .A1(N6207), .B0(N6183));
AND2XL inst_cellmath__34_0_I1978 (.Y(N6236), .A(N6203), .B(N6230));
AOI21XL inst_cellmath__34_0_I1979 (.Y(N6231), .A0(N6263), .A1(N6188), .B0(N6257));
AOI21XL inst_cellmath__34_0_I1980 (.Y(N6245), .A0(N6210), .A1(N6230), .B0(N6207));
AOI31X1 inst_cellmath__34_0_I4144 (.Y(N6177), .A0(N6215), .A1(N6229), .A2(N6178), .B0(N6244));
AOI31X1 inst_cellmath__34_0_I4145 (.Y(N6200), .A0(N6251), .A1(N6261), .A2(N6222), .B0(N6198));
AO21XL inst_cellmath__34_0_I1983 (.Y(N6211), .A0(N6199), .A1(N6263), .B0(N6175));
AO21XL inst_cellmath__34_0_I1984 (.Y(inst_cellmath__34[9]), .A0(N6236), .A1(N6210), .B0(N6220));
NAND2BXL inst_cellmath__34_0_I1985 (.Y(N6197), .AN(N6176), .B(N6254));
NAND2BXL inst_cellmath__34_0_I1986 (.Y(N6252), .AN(N6184), .B(N6204));
NAND2BXL inst_cellmath__34_0_I1987 (.Y(N6226), .AN(N6227), .B(N6240));
NAND2BXL inst_cellmath__34_0_I1988 (.Y(N6192), .AN(N6259), .B(N6193));
NAND2BXL inst_cellmath__34_0_I1989 (.Y(N6248), .AN(N6213), .B(N6232));
NAND2BXL inst_cellmath__34_0_I1990 (.Y(N6223), .AN(N6249), .B(N6180));
NAND2BXL inst_cellmath__34_0_I1991 (.Y(N6190), .AN(N6201), .B(N6224));
XNOR2X1 inst_cellmath__34_0_I1992 (.Y(inst_cellmath__34[0]), .A(N6263), .B(N6218));
XOR2XL inst_cellmath__34_0_I1993 (.Y(inst_cellmath__34[1]), .A(N6210), .B(N6197));
XOR2XL inst_cellmath__34_0_I1994 (.Y(inst_cellmath__34[2]), .A(N6178), .B(N6252));
XOR2XL inst_cellmath__34_0_I1995 (.Y(inst_cellmath__34[3]), .A(N6222), .B(N6226));
XNOR2X1 inst_cellmath__34_0_I1996 (.Y(inst_cellmath__34[4]), .A(N6231), .B(N6192));
XNOR2X1 inst_cellmath__34_0_I1997 (.Y(inst_cellmath__34[5]), .A(N6245), .B(N6248));
XNOR2X1 inst_cellmath__34_0_I1998 (.Y(inst_cellmath__34[6]), .A(N6177), .B(N6223));
XNOR2X1 inst_cellmath__34_0_I1999 (.Y(inst_cellmath__34[7]), .A(N6200), .B(N6190));
XNOR2X1 inst_cellmath__34_0_I2000 (.Y(inst_cellmath__34[8]), .A(N6211), .B(N6189));
AND3XL inst_cellmath__41__24__I4146 (.Y(N6337), .A(inst_cellmath__34[0]), .B(inst_cellmath__34[1]), .C(inst_cellmath__34[2]));
NAND3XL inst_cellmath__41__24__I2003 (.Y(N6349), .A(inst_cellmath__34[3]), .B(N6337), .C(inst_cellmath__34[6]));
NAND3XL inst_cellmath__41__24__I2004 (.Y(N6342), .A(inst_cellmath__34[4]), .B(inst_cellmath__34[7]), .C(inst_cellmath__34[5]));
NOR2XL andori2bb1_A_I4234 (.Y(N9410), .A(N6349), .B(N6342));
NOR2XL andori2bb1_A_I4235 (.Y(N6355), .A(N9410), .B(inst_cellmath__34[8]));
NOR2XL cynw_cm_float_mul_I2009 (.Y(inst_cellmath__41), .A(inst_cellmath__34[9]), .B(N6355));
OR2XL cynw_cm_float_mul_I2010 (.Y(N6367), .A(N6169), .B(inst_cellmath__41));
NOR2XL inst_cellmath__35__16__I2013 (.Y(N6381), .A(inst_cellmath__34[9]), .B(inst_cellmath__34[3]));
NOR2XL inst_cellmath__35__16__I2014 (.Y(N6386), .A(inst_cellmath__34[4]), .B(inst_cellmath__34[6]));
NOR2XL inst_cellmath__35__16__I2015 (.Y(N6389), .A(inst_cellmath__34[5]), .B(inst_cellmath__34[7]));
NOR4X1 inst_cellmath__35__16__I4148 (.Y(N6374), .A(inst_cellmath__34[0]), .B(inst_cellmath__34[1]), .C(inst_cellmath__34[2]), .D(inst_cellmath__34[8]));
NAND4XL inst_cellmath__35__16__I4184 (.Y(N273), .A(N6381), .B(N6389), .C(N6386), .D(N6374));
NOR3BXL cynw_cm_float_mul_I4151 (.Y(N269), .AN(inst_cellmath__25), .B(inst_cellmath__22), .C(inst_cellmath__24));
NOR3BXL cynw_cm_float_mul_I4153 (.Y(N270), .AN(inst_cellmath__26), .B(inst_cellmath__21), .C(inst_cellmath__23));
OR2XL cynw_cm_float_mul_I2026 (.Y(N6417), .A(N269), .B(N270));
NOR3XL inst_cellmath__60_0_I2028 (.Y(N6424), .A(N6417), .B(inst_cellmath__29), .C(inst_cellmath__34[9]));
NAND2XL hyperpropagate_3_1_A_I4236 (.Y(N9417), .A(N6424), .B(N273));
NOR2XL hyperpropagate_3_1_A_I4237 (.Y(N6426), .A(N6367), .B(N9417));
INVXL inst_cellmath__42__22__I2035 (.Y(N6439), .A(inst_cellmath__34[5]));
AND4XL inst_cellmath__42__22__I11248 (.Y(N6437), .A(inst_cellmath__34[3]), .B(inst_cellmath__34[4]), .C(inst_cellmath__34[6]), .D(inst_cellmath__34[7]));
NAND3XL hyperpropagate_4_1_A_I4238 (.Y(N9426), .A(inst_cellmath__34[1]), .B(inst_cellmath__34[2]), .C(N6437));
NOR2XL hyperpropagate_4_1_A_I4239 (.Y(N274), .A(N6439), .B(N9426));
NOR2XL cynw_cm_float_mul_I2039 (.Y(N6457), .A(inst_cellmath__34[8]), .B(N274));
NOR2XL cynw_cm_float_mul_I2042 (.Y(inst_cellmath__42), .A(inst_cellmath__34[9]), .B(N6457));
OR2XL cynw_cm_float_mul_I2043 (.Y(N6469), .A(N6169), .B(inst_cellmath__42));
NOR4X2 cynw_cm_float_mul_I4156 (.Y(N6480), .A(N6469), .B(inst_cellmath__29), .C(inst_cellmath__34[9]), .D(N6417));
INVXL inst_cellmath__50_0_I2052 (.Y(inst_cellmath__50[0]), .A(inst_cellmath__34[0]));
NOR2BX1 inst_cellmath__50_0_I4157 (.Y(N6524), .AN(inst_cellmath__34[1]), .B(inst_cellmath__50[0]));
XNOR2X1 inst_cellmath__50_0_I2054 (.Y(inst_cellmath__50[1]), .A(inst_cellmath__50[0]), .B(inst_cellmath__34[1]));
NAND2XL inst_cellmath__50_0_I2055 (.Y(N6494), .A(inst_cellmath__34[2]), .B(N6524));
NAND2XL inst_cellmath__50_0_I2057 (.Y(N6505), .A(inst_cellmath__34[4]), .B(inst_cellmath__34[3]));
INVXL inst_cellmath__50_0_I2060 (.Y(N6508), .A(N6494));
NOR2XL inst_cellmath__50_0_I2061 (.Y(N6504), .A(N6505), .B(N6494));
NOR4BBX1 inst_cellmath__50_0_I4158 (.Y(N6525), .AN(inst_cellmath__34[6]), .BN(inst_cellmath__34[5]), .C(N6494), .D(N6505));
XOR2XL inst_cellmath__50_0_I2065 (.Y(inst_cellmath__50[2]), .A(N6524), .B(inst_cellmath__34[2]));
XOR2XL inst_cellmath__50_0_I2066 (.Y(inst_cellmath__50[3]), .A(N6508), .B(inst_cellmath__34[3]));
XNOR2X1 inst_cellmath__50_0_I2067 (.Y(inst_cellmath__50[5]), .A(N6504), .B(N6439));
XOR2XL inst_cellmath__50_0_I2068 (.Y(inst_cellmath__50[7]), .A(N6525), .B(inst_cellmath__34[7]));
XOR2XL inst_cellmath__50_0_I4159 (.Y(N6513), .A(inst_cellmath__34[4]), .B(inst_cellmath__34[3]));
MX2XL inst_cellmath__50_0_I4160 (.Y(inst_cellmath__50[4]), .A(inst_cellmath__34[4]), .B(N6513), .S0(N6508));
NAND2BXL inst_cellmath__50_0_I2073 (.Y(N6503), .AN(N6439), .B(N6504));
XNOR2X1 inst_cellmath__50_0_I2074 (.Y(inst_cellmath__50[6]), .A(inst_cellmath__34[6]), .B(N6503));
NOR3XL cynw_cm_float_mul_I2075 (.Y(N6551), .A(inst_cellmath__29), .B(N6367), .C(N6469));
INVXL inst_cellmath__64_2WWMM_I2081 (.Y(N6639), .A(inst_cellmath__29));
INVX2 inst_cellmath__64_2WWMM_I2082 (.Y(N6669), .A(inst_cellmath__43[47]));
CLKINVX4 inst_cellmath__64_2WWMM_I2083 (.Y(N6583), .A(N6669));
MXI2XL inst_cellmath__64_2WWMM_I2089 (.Y(N6652), .A(inst_cellmath__50[0]), .B(inst_cellmath__34[0]), .S0(N6669));
MXI2XL inst_cellmath__64_2WWMM_I2090 (.Y(N6680), .A(inst_cellmath__34[1]), .B(inst_cellmath__50[1]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2091 (.Y(N6581), .A(inst_cellmath__34[2]), .B(inst_cellmath__50[2]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2092 (.Y(N6608), .A(inst_cellmath__34[3]), .B(inst_cellmath__50[3]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2093 (.Y(N6633), .A(inst_cellmath__34[4]), .B(inst_cellmath__50[4]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2094 (.Y(N6663), .A(inst_cellmath__34[5]), .B(inst_cellmath__50[5]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2095 (.Y(N6564), .A(inst_cellmath__34[6]), .B(inst_cellmath__50[6]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2096 (.Y(N6593), .A(inst_cellmath__34[7]), .B(inst_cellmath__50[7]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2097 (.Y(N6618), .A(inst_cellmath__43[23]), .B(inst_cellmath__43[24]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2098 (.Y(N6647), .A(inst_cellmath__43[24]), .B(inst_cellmath__43[25]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2099 (.Y(N6675), .A(inst_cellmath__43[25]), .B(inst_cellmath__43[26]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2100 (.Y(N6575), .A(inst_cellmath__43[26]), .B(inst_cellmath__43[27]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2101 (.Y(N6604), .A(inst_cellmath__43[27]), .B(inst_cellmath__43[28]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2102 (.Y(N6629), .A(inst_cellmath__43[28]), .B(inst_cellmath__43[29]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2103 (.Y(N6659), .A(inst_cellmath__43[29]), .B(inst_cellmath__43[30]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2104 (.Y(N6687), .A(inst_cellmath__43[30]), .B(inst_cellmath__43[31]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2105 (.Y(N6588), .A(inst_cellmath__43[31]), .B(inst_cellmath__43[32]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2106 (.Y(N6613), .A(inst_cellmath__43[32]), .B(inst_cellmath__43[33]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2107 (.Y(N6640), .A(inst_cellmath__43[33]), .B(inst_cellmath__43[34]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2108 (.Y(N6670), .A(inst_cellmath__43[34]), .B(inst_cellmath__43[35]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2109 (.Y(N6571), .A(inst_cellmath__43[35]), .B(inst_cellmath__43[36]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2110 (.Y(N6600), .A(inst_cellmath__43[36]), .B(inst_cellmath__43[37]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2111 (.Y(N6625), .A(inst_cellmath__43[37]), .B(inst_cellmath__43[38]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2112 (.Y(N6654), .A(inst_cellmath__43[38]), .B(inst_cellmath__43[39]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2113 (.Y(N6683), .A(inst_cellmath__43[39]), .B(inst_cellmath__43[40]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2114 (.Y(N6584), .A(inst_cellmath__43[40]), .B(inst_cellmath__43[41]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2115 (.Y(N6610), .A(inst_cellmath__43[41]), .B(inst_cellmath__43[42]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2116 (.Y(N6636), .A(inst_cellmath__43[42]), .B(inst_cellmath__43[43]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2117 (.Y(N6666), .A(inst_cellmath__43[43]), .B(inst_cellmath__43[44]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2118 (.Y(N6567), .A(inst_cellmath__43[44]), .B(inst_cellmath__43[45]), .S0(N6583));
MXI2XL inst_cellmath__64_2WWMM_I2119 (.Y(N6596), .A(inst_cellmath__43[45]), .B(inst_cellmath__43[46]), .S0(N6583));
MXI2X1 inst_cellmath__64_2WWMM_I4076 (.Y(N9354), .A(N6426), .B(N6480), .S0(inst_cellmath__43[47]));
CLKINVX2 inst_cellmath__64_2WWMM_I4065 (.Y(N6635), .A(N9354));
CLKINVX12 inst_cellmath__64_2WWMM_I2121 (.Y(N6578), .A(N6635));
MXI2XL inst_cellmath__64_2WWMM_I2128 (.Y(x[23]), .A(N6652), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2129 (.Y(x[24]), .A(N6680), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2130 (.Y(x[25]), .A(N6581), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2131 (.Y(x[26]), .A(N6608), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2132 (.Y(x[27]), .A(N6633), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2133 (.Y(x[28]), .A(N6663), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2134 (.Y(x[29]), .A(N6564), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2135 (.Y(x[30]), .A(N6593), .B(N6551), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2136 (.Y(x[0]), .A(N6618), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2137 (.Y(x[1]), .A(N6647), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2138 (.Y(x[2]), .A(N6675), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2139 (.Y(x[3]), .A(N6575), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2140 (.Y(x[4]), .A(N6604), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2141 (.Y(x[5]), .A(N6629), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2142 (.Y(x[6]), .A(N6659), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2143 (.Y(x[7]), .A(N6687), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2144 (.Y(x[8]), .A(N6588), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2145 (.Y(x[9]), .A(N6613), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2146 (.Y(x[10]), .A(N6640), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2147 (.Y(x[11]), .A(N6670), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2148 (.Y(x[12]), .A(N6571), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2149 (.Y(x[13]), .A(N6600), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2150 (.Y(x[14]), .A(N6625), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2151 (.Y(x[15]), .A(N6654), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2152 (.Y(x[16]), .A(N6683), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2153 (.Y(x[17]), .A(N6584), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2154 (.Y(x[18]), .A(N6610), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2155 (.Y(x[19]), .A(N6636), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2156 (.Y(x[20]), .A(N6666), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2157 (.Y(x[21]), .A(N6567), .B(N6639), .S0(N6578));
MXI2XL inst_cellmath__64_2WWMM_I2158 (.Y(x[22]), .A(N6596), .B(N6639), .S0(N6578));
assign inst_cellmath__43[0] = 1'B0;
assign inst_cellmath__43[1] = 1'B0;
assign inst_cellmath__43[2] = 1'B0;
assign inst_cellmath__43[3] = 1'B0;
assign inst_cellmath__43[4] = 1'B0;
assign inst_cellmath__43[5] = 1'B0;
assign inst_cellmath__43[6] = 1'B0;
assign inst_cellmath__43[7] = 1'B0;
assign inst_cellmath__43[8] = 1'B0;
assign inst_cellmath__43[9] = 1'B0;
assign inst_cellmath__43[10] = 1'B0;
assign inst_cellmath__43[11] = 1'B0;
assign inst_cellmath__43[12] = 1'B0;
assign inst_cellmath__43[13] = 1'B0;
assign inst_cellmath__43[14] = 1'B0;
assign inst_cellmath__43[15] = 1'B0;
assign inst_cellmath__43[16] = 1'B0;
assign inst_cellmath__43[17] = 1'B0;
assign inst_cellmath__43[18] = 1'B0;
assign inst_cellmath__43[19] = 1'B0;
assign inst_cellmath__43[20] = 1'B0;
assign inst_cellmath__43[21] = 1'B0;
assign inst_cellmath__43[22] = 1'B0;
endmodule

/* CADENCE  urfwSA/Zoxw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



